// DE4_SOPC.v

// Generated using ACDS version 12.1 177 at 2013.01.18.12:06:11

`timescale 1 ps / 1 ps
module DE4_SOPC (
		output wire        sram_clk_clk,                    //                 sram_clk.clk
		input  wire [15:0] switches_export,                 //                 switches.export
		input  wire        clk_50,                          //            clk_50_clk_in.clk
		input  wire [9:0]  touch_x1,                        //                    touch.x1
		input  wire [8:0]  touch_y1,                        //                         .y1
		input  wire [9:0]  touch_x2,                        //                         .x2
		input  wire [8:0]  touch_y2,                        //                         .y2
		input  wire [9:0]  touch_count_gesture,             //                         .count_gesture
		input  wire        touch_touch_valid,               //                         .touch_valid
		output wire        mem_ssram_adv,                   //                      mem.ssram_adv
		output wire        mem_ssram_bwa_n,                 //                         .ssram_bwa_n
		output wire        mem_ssram_bwb_n,                 //                         .ssram_bwb_n
		output wire        mem_ssram_ce_n,                  //                         .ssram_ce_n
		output wire        mem_ssram_cke_n,                 //                         .ssram_cke_n
		output wire        mem_ssram_oe_n,                  //                         .ssram_oe_n
		output wire        mem_ssram_we_n,                  //                         .ssram_we_n
		output wire [24:0] mem_fsm_a,                       //                         .fsm_a
		output wire [15:0] mem_fsm_d_out,                   //                         .fsm_d_out
		input  wire [15:0] mem_fsm_d_in,                    //                         .fsm_d_in
		output wire        mem_fsm_dout_req,                //                         .fsm_dout_req
		output wire        mem_flash_adv_n,                 //                         .flash_adv_n
		output wire        mem_flash_ce_n,                  //                         .flash_ce_n
		output wire        mem_flash_clk,                   //                         .flash_clk
		output wire        mem_flash_oe_n,                  //                         .flash_oe_n
		output wire        mem_flash_we_n,                  //                         .flash_we_n
		inout  wire        sd_b_SD_cmd,                     //                       sd.b_SD_cmd
		inout  wire        sd_b_SD_dat,                     //                         .b_SD_dat
		inout  wire        sd_b_SD_dat3,                    //                         .b_SD_dat3
		output wire        sd_o_SD_clock,                   //                         .o_SD_clock
		input  wire        reset_reset_n,                   //                    reset.reset_n
		output wire [7:0]  leds_external_connection_export, // leds_external_connection.export
		output wire [7:0]  mtl_lcd_r,                       //                  mtl_lcd.r
		output wire [7:0]  mtl_lcd_g,                       //                         .g
		output wire [7:0]  mtl_lcd_b,                       //                         .b
		output wire        mtl_lcd_hsd,                     //                         .hsd
		output wire        mtl_lcd_vsd                      //                         .vsd
	);

	wire          timing_adapter_1_out_endofpacket;                                                                                         // timing_adapter_1:out_endofpacket -> receive_fifo:avalonst_sink_endofpacket
	wire          timing_adapter_1_out_valid;                                                                                               // timing_adapter_1:out_valid -> receive_fifo:avalonst_sink_valid
	wire          timing_adapter_1_out_startofpacket;                                                                                       // timing_adapter_1:out_startofpacket -> receive_fifo:avalonst_sink_startofpacket
	wire    [5:0] timing_adapter_1_out_error;                                                                                               // timing_adapter_1:out_error -> receive_fifo:avalonst_sink_error
	wire    [1:0] timing_adapter_1_out_empty;                                                                                               // timing_adapter_1:out_empty -> receive_fifo:avalonst_sink_empty
	wire   [31:0] timing_adapter_1_out_data;                                                                                                // timing_adapter_1:out_data -> receive_fifo:avalonst_sink_data
	wire          timing_adapter_1_out_ready;                                                                                               // receive_fifo:avalonst_sink_ready -> timing_adapter_1:out_ready
	wire          dc_fifo_0_out_endofpacket;                                                                                                // dc_fifo_0:out_endofpacket -> AvalonStream2MTL_LCD24bit_0:asi_stream_in_endofpacket
	wire          dc_fifo_0_out_valid;                                                                                                      // dc_fifo_0:out_valid -> AvalonStream2MTL_LCD24bit_0:asi_stream_in_valid
	wire          dc_fifo_0_out_startofpacket;                                                                                              // dc_fifo_0:out_startofpacket -> AvalonStream2MTL_LCD24bit_0:asi_stream_in_startofpacket
	wire   [23:0] dc_fifo_0_out_data;                                                                                                       // dc_fifo_0:out_data -> AvalonStream2MTL_LCD24bit_0:asi_stream_in_data
	wire          dc_fifo_0_out_ready;                                                                                                      // AvalonStream2MTL_LCD24bit_0:asi_stream_in_ready -> dc_fifo_0:out_ready
	wire          mkmtl_framebuffer_flash_0_stream_out_endofpacket;                                                                         // mkMTL_Framebuffer_Flash_0:aso_stream_out_endofpacket -> dc_fifo_0:in_endofpacket
	wire          mkmtl_framebuffer_flash_0_stream_out_valid;                                                                               // mkMTL_Framebuffer_Flash_0:aso_stream_out_valid -> dc_fifo_0:in_valid
	wire          mkmtl_framebuffer_flash_0_stream_out_startofpacket;                                                                       // mkMTL_Framebuffer_Flash_0:aso_stream_out_startofpacket -> dc_fifo_0:in_startofpacket
	wire   [23:0] mkmtl_framebuffer_flash_0_stream_out_data;                                                                                // mkMTL_Framebuffer_Flash_0:aso_stream_out_data -> dc_fifo_0:in_data
	wire          mkmtl_framebuffer_flash_0_stream_out_ready;                                                                               // dc_fifo_0:in_ready -> mkMTL_Framebuffer_Flash_0:aso_stream_out_ready
	wire          transmit_fifo_out_endofpacket;                                                                                            // transmit_fifo:avalonst_source_endofpacket -> timing_adapter:in_endofpacket
	wire          transmit_fifo_out_valid;                                                                                                  // transmit_fifo:avalonst_source_valid -> timing_adapter:in_valid
	wire          transmit_fifo_out_startofpacket;                                                                                          // transmit_fifo:avalonst_source_startofpacket -> timing_adapter:in_startofpacket
	wire          transmit_fifo_out_error;                                                                                                  // transmit_fifo:avalonst_source_error -> timing_adapter:in_error
	wire    [1:0] transmit_fifo_out_empty;                                                                                                  // transmit_fifo:avalonst_source_empty -> timing_adapter:in_empty
	wire   [31:0] transmit_fifo_out_data;                                                                                                   // transmit_fifo:avalonst_source_data -> timing_adapter:in_data
	wire          transmit_fifo_out_ready;                                                                                                  // timing_adapter:in_ready -> transmit_fifo:avalonst_source_ready
	wire    [0:0] peripheral_bridge_m0_burstcount;                                                                                          // peripheral_bridge:m0_burstcount -> peripheral_bridge_m0_translator:av_burstcount
	wire          peripheral_bridge_m0_waitrequest;                                                                                         // peripheral_bridge_m0_translator:av_waitrequest -> peripheral_bridge:m0_waitrequest
	wire   [29:0] peripheral_bridge_m0_address;                                                                                             // peripheral_bridge:m0_address -> peripheral_bridge_m0_translator:av_address
	wire   [31:0] peripheral_bridge_m0_writedata;                                                                                           // peripheral_bridge:m0_writedata -> peripheral_bridge_m0_translator:av_writedata
	wire          peripheral_bridge_m0_write;                                                                                               // peripheral_bridge:m0_write -> peripheral_bridge_m0_translator:av_write
	wire          peripheral_bridge_m0_read;                                                                                                // peripheral_bridge:m0_read -> peripheral_bridge_m0_translator:av_read
	wire   [31:0] peripheral_bridge_m0_readdata;                                                                                            // peripheral_bridge_m0_translator:av_readdata -> peripheral_bridge:m0_readdata
	wire          peripheral_bridge_m0_debugaccess;                                                                                         // peripheral_bridge:m0_debugaccess -> peripheral_bridge_m0_translator:av_debugaccess
	wire    [3:0] peripheral_bridge_m0_byteenable;                                                                                          // peripheral_bridge:m0_byteenable -> peripheral_bridge_m0_translator:av_byteenable
	wire          peripheral_bridge_m0_readdatavalid;                                                                                       // peripheral_bridge_m0_translator:av_readdatavalid -> peripheral_bridge:m0_readdatavalid
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_waitrequest;                                                 // mm_clock_crossing_bridge_0:s0_waitrequest -> mm_clock_crossing_bridge_0_s0_translator:av_waitrequest
	wire    [0:0] mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_burstcount;                                                  // mm_clock_crossing_bridge_0_s0_translator:av_burstcount -> mm_clock_crossing_bridge_0:s0_burstcount
	wire   [31:0] mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_writedata;                                                   // mm_clock_crossing_bridge_0_s0_translator:av_writedata -> mm_clock_crossing_bridge_0:s0_writedata
	wire   [17:0] mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_address;                                                     // mm_clock_crossing_bridge_0_s0_translator:av_address -> mm_clock_crossing_bridge_0:s0_address
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_write;                                                       // mm_clock_crossing_bridge_0_s0_translator:av_write -> mm_clock_crossing_bridge_0:s0_write
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_read;                                                        // mm_clock_crossing_bridge_0_s0_translator:av_read -> mm_clock_crossing_bridge_0:s0_read
	wire   [31:0] mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdata;                                                    // mm_clock_crossing_bridge_0:s0_readdata -> mm_clock_crossing_bridge_0_s0_translator:av_readdata
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_debugaccess;                                                 // mm_clock_crossing_bridge_0_s0_translator:av_debugaccess -> mm_clock_crossing_bridge_0:s0_debugaccess
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdatavalid;                                               // mm_clock_crossing_bridge_0:s0_readdatavalid -> mm_clock_crossing_bridge_0_s0_translator:av_readdatavalid
	wire    [3:0] mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_byteenable;                                                  // mm_clock_crossing_bridge_0_s0_translator:av_byteenable -> mm_clock_crossing_bridge_0:s0_byteenable
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_waitrequest;                                                  // mkMTL_Framebuffer_Flash_0:avs_s0_waitrequest -> mkMTL_Framebuffer_Flash_0_s0_translator:av_waitrequest
	wire   [31:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_writedata;                                                    // mkMTL_Framebuffer_Flash_0_s0_translator:av_writedata -> mkMTL_Framebuffer_Flash_0:avs_s0_writedata
	wire   [24:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_address;                                                      // mkMTL_Framebuffer_Flash_0_s0_translator:av_address -> mkMTL_Framebuffer_Flash_0:avs_s0_address
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_write;                                                        // mkMTL_Framebuffer_Flash_0_s0_translator:av_write -> mkMTL_Framebuffer_Flash_0:avs_s0_write
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_read;                                                         // mkMTL_Framebuffer_Flash_0_s0_translator:av_read -> mkMTL_Framebuffer_Flash_0:avs_s0_read
	wire   [31:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_readdata;                                                     // mkMTL_Framebuffer_Flash_0:avs_s0_readdata -> mkMTL_Framebuffer_Flash_0_s0_translator:av_readdata
	wire    [3:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_byteenable;                                                   // mkMTL_Framebuffer_Flash_0_s0_translator:av_byteenable -> mkMTL_Framebuffer_Flash_0:avs_s0_byteenable
	wire   [31:0] onchip_memory_mips_s1_translator_avalon_anti_slave_0_writedata;                                                           // onchip_memory_MIPS_s1_translator:av_writedata -> onchip_memory_MIPS:writedata
	wire   [12:0] onchip_memory_mips_s1_translator_avalon_anti_slave_0_address;                                                             // onchip_memory_MIPS_s1_translator:av_address -> onchip_memory_MIPS:address
	wire          onchip_memory_mips_s1_translator_avalon_anti_slave_0_chipselect;                                                          // onchip_memory_MIPS_s1_translator:av_chipselect -> onchip_memory_MIPS:chipselect
	wire          onchip_memory_mips_s1_translator_avalon_anti_slave_0_clken;                                                               // onchip_memory_MIPS_s1_translator:av_clken -> onchip_memory_MIPS:clken
	wire          onchip_memory_mips_s1_translator_avalon_anti_slave_0_write;                                                               // onchip_memory_MIPS_s1_translator:av_write -> onchip_memory_MIPS:write
	wire   [31:0] onchip_memory_mips_s1_translator_avalon_anti_slave_0_readdata;                                                            // onchip_memory_MIPS:readdata -> onchip_memory_MIPS_s1_translator:av_readdata
	wire    [3:0] onchip_memory_mips_s1_translator_avalon_anti_slave_0_byteenable;                                                          // onchip_memory_MIPS_s1_translator:av_byteenable -> onchip_memory_MIPS:byteenable
	wire    [0:0] mm_clock_crossing_bridge_0_m0_burstcount;                                                                                 // mm_clock_crossing_bridge_0:m0_burstcount -> mm_clock_crossing_bridge_0_m0_translator:av_burstcount
	wire          mm_clock_crossing_bridge_0_m0_waitrequest;                                                                                // mm_clock_crossing_bridge_0_m0_translator:av_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	wire   [17:0] mm_clock_crossing_bridge_0_m0_address;                                                                                    // mm_clock_crossing_bridge_0:m0_address -> mm_clock_crossing_bridge_0_m0_translator:av_address
	wire   [31:0] mm_clock_crossing_bridge_0_m0_writedata;                                                                                  // mm_clock_crossing_bridge_0:m0_writedata -> mm_clock_crossing_bridge_0_m0_translator:av_writedata
	wire          mm_clock_crossing_bridge_0_m0_write;                                                                                      // mm_clock_crossing_bridge_0:m0_write -> mm_clock_crossing_bridge_0_m0_translator:av_write
	wire          mm_clock_crossing_bridge_0_m0_read;                                                                                       // mm_clock_crossing_bridge_0:m0_read -> mm_clock_crossing_bridge_0_m0_translator:av_read
	wire   [31:0] mm_clock_crossing_bridge_0_m0_readdata;                                                                                   // mm_clock_crossing_bridge_0_m0_translator:av_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	wire          mm_clock_crossing_bridge_0_m0_debugaccess;                                                                                // mm_clock_crossing_bridge_0:m0_debugaccess -> mm_clock_crossing_bridge_0_m0_translator:av_debugaccess
	wire    [3:0] mm_clock_crossing_bridge_0_m0_byteenable;                                                                                 // mm_clock_crossing_bridge_0:m0_byteenable -> mm_clock_crossing_bridge_0_m0_translator:av_byteenable
	wire          mm_clock_crossing_bridge_0_m0_readdatavalid;                                                                              // mm_clock_crossing_bridge_0_m0_translator:av_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest;                           // Altera_UP_SD_Card_Avalon_Interface_1:o_avalon_waitrequest -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:av_waitrequest
	wire   [31:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                             // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:av_writedata -> Altera_UP_SD_Card_Avalon_Interface_1:i_avalon_writedata
	wire    [7:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_address;                               // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:av_address -> Altera_UP_SD_Card_Avalon_Interface_1:i_avalon_address
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                            // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:av_chipselect -> Altera_UP_SD_Card_Avalon_Interface_1:i_avalon_chip_select
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_write;                                 // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:av_write -> Altera_UP_SD_Card_Avalon_Interface_1:i_avalon_write
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_read;                                  // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:av_read -> Altera_UP_SD_Card_Avalon_Interface_1:i_avalon_read
	wire   [31:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                              // Altera_UP_SD_Card_Avalon_Interface_1:o_avalon_readdata -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:av_readdata
	wire    [3:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                            // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:av_byteenable -> Altera_UP_SD_Card_Avalon_Interface_1:i_avalon_byteenable
	wire   [31:0] leds_s1_translator_avalon_anti_slave_0_writedata;                                                                         // LEDs_s1_translator:av_writedata -> LEDs:writedata
	wire    [1:0] leds_s1_translator_avalon_anti_slave_0_address;                                                                           // LEDs_s1_translator:av_address -> LEDs:address
	wire          leds_s1_translator_avalon_anti_slave_0_chipselect;                                                                        // LEDs_s1_translator:av_chipselect -> LEDs:chipselect
	wire          leds_s1_translator_avalon_anti_slave_0_write;                                                                             // LEDs_s1_translator:av_write -> LEDs:write_n
	wire   [31:0] leds_s1_translator_avalon_anti_slave_0_readdata;                                                                          // LEDs:readdata -> LEDs_s1_translator:av_readdata
	wire    [1:0] switches_s1_translator_avalon_anti_slave_0_address;                                                                       // Switches_s1_translator:av_address -> Switches:address
	wire   [31:0] switches_s1_translator_avalon_anti_slave_0_readdata;                                                                      // Switches:readdata -> Switches_s1_translator:av_readdata
	wire          transmit_fifo_in_translator_avalon_anti_slave_0_waitrequest;                                                              // transmit_fifo:avalonmm_write_slave_waitrequest -> transmit_fifo_in_translator:av_waitrequest
	wire   [31:0] transmit_fifo_in_translator_avalon_anti_slave_0_writedata;                                                                // transmit_fifo_in_translator:av_writedata -> transmit_fifo:avalonmm_write_slave_writedata
	wire    [0:0] transmit_fifo_in_translator_avalon_anti_slave_0_address;                                                                  // transmit_fifo_in_translator:av_address -> transmit_fifo:avalonmm_write_slave_address
	wire          transmit_fifo_in_translator_avalon_anti_slave_0_write;                                                                    // transmit_fifo_in_translator:av_write -> transmit_fifo:avalonmm_write_slave_write
	wire   [31:0] transmit_fifo_in_csr_translator_avalon_anti_slave_0_writedata;                                                            // transmit_fifo_in_csr_translator:av_writedata -> transmit_fifo:wrclk_control_slave_writedata
	wire    [2:0] transmit_fifo_in_csr_translator_avalon_anti_slave_0_address;                                                              // transmit_fifo_in_csr_translator:av_address -> transmit_fifo:wrclk_control_slave_address
	wire          transmit_fifo_in_csr_translator_avalon_anti_slave_0_write;                                                                // transmit_fifo_in_csr_translator:av_write -> transmit_fifo:wrclk_control_slave_write
	wire          transmit_fifo_in_csr_translator_avalon_anti_slave_0_read;                                                                 // transmit_fifo_in_csr_translator:av_read -> transmit_fifo:wrclk_control_slave_read
	wire   [31:0] transmit_fifo_in_csr_translator_avalon_anti_slave_0_readdata;                                                             // transmit_fifo:wrclk_control_slave_readdata -> transmit_fifo_in_csr_translator:av_readdata
	wire          receive_fifo_out_translator_avalon_anti_slave_0_waitrequest;                                                              // receive_fifo:avalonmm_read_slave_waitrequest -> receive_fifo_out_translator:av_waitrequest
	wire    [0:0] receive_fifo_out_translator_avalon_anti_slave_0_address;                                                                  // receive_fifo_out_translator:av_address -> receive_fifo:avalonmm_read_slave_address
	wire          receive_fifo_out_translator_avalon_anti_slave_0_read;                                                                     // receive_fifo_out_translator:av_read -> receive_fifo:avalonmm_read_slave_read
	wire   [31:0] receive_fifo_out_translator_avalon_anti_slave_0_readdata;                                                                 // receive_fifo:avalonmm_read_slave_readdata -> receive_fifo_out_translator:av_readdata
	wire   [31:0] receive_fifo_out_csr_translator_avalon_anti_slave_0_writedata;                                                            // receive_fifo_out_csr_translator:av_writedata -> receive_fifo:rdclk_control_slave_writedata
	wire    [2:0] receive_fifo_out_csr_translator_avalon_anti_slave_0_address;                                                              // receive_fifo_out_csr_translator:av_address -> receive_fifo:rdclk_control_slave_address
	wire          receive_fifo_out_csr_translator_avalon_anti_slave_0_write;                                                                // receive_fifo_out_csr_translator:av_write -> receive_fifo:rdclk_control_slave_write
	wire          receive_fifo_out_csr_translator_avalon_anti_slave_0_read;                                                                 // receive_fifo_out_csr_translator:av_read -> receive_fifo:rdclk_control_slave_read
	wire   [31:0] receive_fifo_out_csr_translator_avalon_anti_slave_0_readdata;                                                             // receive_fifo:rdclk_control_slave_readdata -> receive_fifo_out_csr_translator:av_readdata
	wire   [31:0] versionrom_s1_translator_avalon_anti_slave_0_writedata;                                                                   // versionRom_s1_translator:av_writedata -> versionRom:writedata
	wire    [2:0] versionrom_s1_translator_avalon_anti_slave_0_address;                                                                     // versionRom_s1_translator:av_address -> versionRom:address
	wire          versionrom_s1_translator_avalon_anti_slave_0_chipselect;                                                                  // versionRom_s1_translator:av_chipselect -> versionRom:chipselect
	wire          versionrom_s1_translator_avalon_anti_slave_0_clken;                                                                       // versionRom_s1_translator:av_clken -> versionRom:clken
	wire          versionrom_s1_translator_avalon_anti_slave_0_write;                                                                       // versionRom_s1_translator:av_write -> versionRom:write
	wire   [31:0] versionrom_s1_translator_avalon_anti_slave_0_readdata;                                                                    // versionRom:readdata -> versionRom_s1_translator:av_readdata
	wire          versionrom_s1_translator_avalon_anti_slave_0_debugaccess;                                                                 // versionRom_s1_translator:av_debugaccess -> versionRom:debugaccess
	wire    [3:0] versionrom_s1_translator_avalon_anti_slave_0_byteenable;                                                                  // versionRom_s1_translator:av_byteenable -> versionRom:byteenable
	wire          cheri_avalon_master_0_waitrequest;                                                                                        // CHERI_avalon_master_0_translator:av_waitrequest -> CHERI:avm_waitrequest
	wire   [31:0] cheri_avalon_master_0_address;                                                                                            // CHERI:avm_address -> CHERI_avalon_master_0_translator:av_address
	wire  [255:0] cheri_avalon_master_0_writedata;                                                                                          // CHERI:avm_writedata -> CHERI_avalon_master_0_translator:av_writedata
	wire          cheri_avalon_master_0_write;                                                                                              // CHERI:avm_write -> CHERI_avalon_master_0_translator:av_write
	wire          cheri_avalon_master_0_read;                                                                                               // CHERI:avm_read -> CHERI_avalon_master_0_translator:av_read
	wire  [255:0] cheri_avalon_master_0_readdata;                                                                                           // CHERI_avalon_master_0_translator:av_readdata -> CHERI:avm_readdata
	wire   [31:0] cheri_avalon_master_0_byteenable;                                                                                         // CHERI:avm_byteenable -> CHERI_avalon_master_0_translator:av_byteenable
	wire          cheri_avalon_master_0_readdatavalid;                                                                                      // CHERI_avalon_master_0_translator:av_readdatavalid -> CHERI:avm_readdatavalid
	wire          peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                                          // peripheral_bridge:s0_waitrequest -> peripheral_bridge_s0_translator:av_waitrequest
	wire    [0:0] peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                                           // peripheral_bridge_s0_translator:av_burstcount -> peripheral_bridge:s0_burstcount
	wire   [31:0] peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata;                                                            // peripheral_bridge_s0_translator:av_writedata -> peripheral_bridge:s0_writedata
	wire   [29:0] peripheral_bridge_s0_translator_avalon_anti_slave_0_address;                                                              // peripheral_bridge_s0_translator:av_address -> peripheral_bridge:s0_address
	wire          peripheral_bridge_s0_translator_avalon_anti_slave_0_write;                                                                // peripheral_bridge_s0_translator:av_write -> peripheral_bridge:s0_write
	wire          peripheral_bridge_s0_translator_avalon_anti_slave_0_read;                                                                 // peripheral_bridge_s0_translator:av_read -> peripheral_bridge:s0_read
	wire   [31:0] peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata;                                                             // peripheral_bridge:s0_readdata -> peripheral_bridge_s0_translator:av_readdata
	wire          peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                                          // peripheral_bridge_s0_translator:av_debugaccess -> peripheral_bridge:s0_debugaccess
	wire          peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                                        // peripheral_bridge:s0_readdatavalid -> peripheral_bridge_s0_translator:av_readdatavalid
	wire    [3:0] peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                                           // peripheral_bridge_s0_translator:av_byteenable -> peripheral_bridge:s0_byteenable
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest;                                                    // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> peripheral_bridge_m0_translator:uav_waitrequest
	wire    [2:0] peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount;                                                     // peripheral_bridge_m0_translator:uav_burstcount -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] peripheral_bridge_m0_translator_avalon_universal_master_0_writedata;                                                      // peripheral_bridge_m0_translator:uav_writedata -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [29:0] peripheral_bridge_m0_translator_avalon_universal_master_0_address;                                                        // peripheral_bridge_m0_translator:uav_address -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_lock;                                                           // peripheral_bridge_m0_translator:uav_lock -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_write;                                                          // peripheral_bridge_m0_translator:uav_write -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_read;                                                           // peripheral_bridge_m0_translator:uav_read -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] peripheral_bridge_m0_translator_avalon_universal_master_0_readdata;                                                       // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> peripheral_bridge_m0_translator:uav_readdata
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess;                                                    // peripheral_bridge_m0_translator:uav_debugaccess -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable;                                                     // peripheral_bridge_m0_translator:uav_byteenable -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                                                  // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> peripheral_bridge_m0_translator:uav_readdatavalid
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // mm_clock_crossing_bridge_0_s0_translator:uav_waitrequest -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> mm_clock_crossing_bridge_0_s0_translator:uav_burstcount
	wire   [31:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> mm_clock_crossing_bridge_0_s0_translator:uav_writedata
	wire   [29:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_address;                                       // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_address -> mm_clock_crossing_bridge_0_s0_translator:uav_address
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_write;                                         // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_write -> mm_clock_crossing_bridge_0_s0_translator:uav_write
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                          // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_lock -> mm_clock_crossing_bridge_0_s0_translator:uav_lock
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_read;                                          // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_read -> mm_clock_crossing_bridge_0_s0_translator:uav_read
	wire   [31:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // mm_clock_crossing_bridge_0_s0_translator:uav_readdata -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // mm_clock_crossing_bridge_0_s0_translator:uav_readdatavalid -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mm_clock_crossing_bridge_0_s0_translator:uav_debugaccess
	wire    [3:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> mm_clock_crossing_bridge_0_s0_translator:uav_byteenable
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // mkMTL_Framebuffer_Flash_0_s0_translator:uav_waitrequest -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> mkMTL_Framebuffer_Flash_0_s0_translator:uav_burstcount
	wire   [31:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> mkMTL_Framebuffer_Flash_0_s0_translator:uav_writedata
	wire   [29:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_address;                                        // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_address -> mkMTL_Framebuffer_Flash_0_s0_translator:uav_address
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_write;                                          // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_write -> mkMTL_Framebuffer_Flash_0_s0_translator:uav_write
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                           // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_lock -> mkMTL_Framebuffer_Flash_0_s0_translator:uav_lock
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_read;                                           // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_read -> mkMTL_Framebuffer_Flash_0_s0_translator:uav_read
	wire   [31:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // mkMTL_Framebuffer_Flash_0_s0_translator:uav_readdata -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // mkMTL_Framebuffer_Flash_0_s0_translator:uav_readdatavalid -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mkMTL_Framebuffer_Flash_0_s0_translator:uav_debugaccess
	wire    [3:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> mkMTL_Framebuffer_Flash_0_s0_translator:uav_byteenable
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                           // onchip_memory_MIPS_s1_translator:uav_waitrequest -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                            // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory_MIPS_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                             // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory_MIPS_s1_translator:uav_writedata
	wire   [29:0] onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_address;                                               // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory_MIPS_s1_translator:uav_address
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                 // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory_MIPS_s1_translator:uav_write
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                  // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory_MIPS_s1_translator:uav_lock
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                  // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory_MIPS_s1_translator:uav_read
	wire   [31:0] onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                              // onchip_memory_MIPS_s1_translator:uav_readdata -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                         // onchip_memory_MIPS_s1_translator:uav_readdatavalid -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                           // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory_MIPS_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                            // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory_MIPS_s1_translator:uav_byteenable
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                    // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                          // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                  // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                           // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                          // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                 // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                       // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                               // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                        // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                       // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                     // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                      // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                     // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_waitrequest;                                           // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> mm_clock_crossing_bridge_0_m0_translator:uav_waitrequest
	wire    [2:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_burstcount;                                            // mm_clock_crossing_bridge_0_m0_translator:uav_burstcount -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_writedata;                                             // mm_clock_crossing_bridge_0_m0_translator:uav_writedata -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [17:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_address;                                               // mm_clock_crossing_bridge_0_m0_translator:uav_address -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_address
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_lock;                                                  // mm_clock_crossing_bridge_0_m0_translator:uav_lock -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_write;                                                 // mm_clock_crossing_bridge_0_m0_translator:uav_write -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_write
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_read;                                                  // mm_clock_crossing_bridge_0_m0_translator:uav_read -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdata;                                              // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_readdata -> mm_clock_crossing_bridge_0_m0_translator:uav_readdata
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_debugaccess;                                           // mm_clock_crossing_bridge_0_m0_translator:uav_debugaccess -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_byteenable;                                            // mm_clock_crossing_bridge_0_m0_translator:uav_byteenable -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdatavalid;                                         // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> mm_clock_crossing_bridge_0_m0_translator:uav_readdatavalid
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_waitrequest -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;               // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_writedata
	wire   [17:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                 // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_address
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                   // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_write
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                    // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_lock
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                    // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_read
	wire   [31:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_readdata -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_readdatavalid -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:uav_byteenable
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;             // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                         // LEDs_s1_translator:uav_waitrequest -> LEDs_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                          // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LEDs_s1_translator:uav_burstcount
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                           // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LEDs_s1_translator:uav_writedata
	wire   [17:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                             // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_address -> LEDs_s1_translator:uav_address
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                               // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_write -> LEDs_s1_translator:uav_write
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LEDs_s1_translator:uav_lock
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_read -> LEDs_s1_translator:uav_read
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                            // LEDs_s1_translator:uav_readdata -> LEDs_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                       // LEDs_s1_translator:uav_readdatavalid -> LEDs_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                         // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LEDs_s1_translator:uav_debugaccess
	wire    [3:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                          // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LEDs_s1_translator:uav_byteenable
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                  // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                        // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                         // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                        // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                               // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                     // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                             // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                      // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                     // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                   // LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                    // LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                   // LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                     // Switches_s1_translator:uav_waitrequest -> Switches_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                      // Switches_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Switches_s1_translator:uav_burstcount
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                       // Switches_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Switches_s1_translator:uav_writedata
	wire   [17:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                         // Switches_s1_translator_avalon_universal_slave_0_agent:m0_address -> Switches_s1_translator:uav_address
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                           // Switches_s1_translator_avalon_universal_slave_0_agent:m0_write -> Switches_s1_translator:uav_write
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                            // Switches_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Switches_s1_translator:uav_lock
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                            // Switches_s1_translator_avalon_universal_slave_0_agent:m0_read -> Switches_s1_translator:uav_read
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                        // Switches_s1_translator:uav_readdata -> Switches_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                   // Switches_s1_translator:uav_readdatavalid -> Switches_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                     // Switches_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Switches_s1_translator:uav_debugaccess
	wire    [3:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                      // Switches_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Switches_s1_translator:uav_byteenable
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                              // Switches_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                    // Switches_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                            // Switches_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                     // Switches_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                    // Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Switches_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                           // Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                 // Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                         // Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                  // Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                 // Switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                               // Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                // Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                               // Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // transmit_fifo_in_translator:uav_waitrequest -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> transmit_fifo_in_translator:uav_burstcount
	wire   [31:0] transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_writedata -> transmit_fifo_in_translator:uav_writedata
	wire   [17:0] transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_address;                                                    // transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_address -> transmit_fifo_in_translator:uav_address
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_write;                                                      // transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_write -> transmit_fifo_in_translator:uav_write
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_lock -> transmit_fifo_in_translator:uav_lock
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_read;                                                       // transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_read -> transmit_fifo_in_translator:uav_read
	wire   [31:0] transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // transmit_fifo_in_translator:uav_readdata -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // transmit_fifo_in_translator:uav_readdatavalid -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> transmit_fifo_in_translator:uav_debugaccess
	wire    [3:0] transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // transmit_fifo_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> transmit_fifo_in_translator:uav_byteenable
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rf_source_data -> transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] transmit_fifo_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                            // transmit_fifo_in_csr_translator:uav_waitrequest -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                                             // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> transmit_fifo_in_csr_translator:uav_burstcount
	wire   [31:0] transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                              // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> transmit_fifo_in_csr_translator:uav_writedata
	wire   [17:0] transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                                // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> transmit_fifo_in_csr_translator:uav_address
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                                  // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> transmit_fifo_in_csr_translator:uav_write
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                                   // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> transmit_fifo_in_csr_translator:uav_lock
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                                   // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> transmit_fifo_in_csr_translator:uav_read
	wire   [31:0] transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                               // transmit_fifo_in_csr_translator:uav_readdata -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                          // transmit_fifo_in_csr_translator:uav_readdatavalid -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                            // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> transmit_fifo_in_csr_translator:uav_debugaccess
	wire    [3:0] transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                                             // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> transmit_fifo_in_csr_translator:uav_byteenable
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                     // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                                           // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                   // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                                            // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                                           // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                  // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                        // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                         // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                        // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                      // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                       // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                      // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // receive_fifo_out_translator:uav_waitrequest -> receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> receive_fifo_out_translator:uav_burstcount
	wire   [31:0] receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_writedata -> receive_fifo_out_translator:uav_writedata
	wire   [17:0] receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_address;                                                    // receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_address -> receive_fifo_out_translator:uav_address
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_write;                                                      // receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_write -> receive_fifo_out_translator:uav_write
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_lock -> receive_fifo_out_translator:uav_lock
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_read;                                                       // receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_read -> receive_fifo_out_translator:uav_read
	wire   [31:0] receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // receive_fifo_out_translator:uav_readdata -> receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // receive_fifo_out_translator:uav_readdatavalid -> receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> receive_fifo_out_translator:uav_debugaccess
	wire    [3:0] receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // receive_fifo_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> receive_fifo_out_translator:uav_byteenable
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // receive_fifo_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // receive_fifo_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // receive_fifo_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // receive_fifo_out_translator_avalon_universal_slave_0_agent:rf_source_data -> receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> receive_fifo_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> receive_fifo_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> receive_fifo_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> receive_fifo_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> receive_fifo_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // receive_fifo_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // receive_fifo_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> receive_fifo_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] receive_fifo_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // receive_fifo_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> receive_fifo_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // receive_fifo_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> receive_fifo_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                            // receive_fifo_out_csr_translator:uav_waitrequest -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                                             // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> receive_fifo_out_csr_translator:uav_burstcount
	wire   [31:0] receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                              // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> receive_fifo_out_csr_translator:uav_writedata
	wire   [17:0] receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_address;                                                // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_address -> receive_fifo_out_csr_translator:uav_address
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_write;                                                  // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_write -> receive_fifo_out_csr_translator:uav_write
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                                   // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_lock -> receive_fifo_out_csr_translator:uav_lock
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_read;                                                   // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_read -> receive_fifo_out_csr_translator:uav_read
	wire   [31:0] receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                               // receive_fifo_out_csr_translator:uav_readdata -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                          // receive_fifo_out_csr_translator:uav_readdatavalid -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                            // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> receive_fifo_out_csr_translator:uav_debugaccess
	wire    [3:0] receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                                             // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> receive_fifo_out_csr_translator:uav_byteenable
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                     // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                                           // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                   // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                                            // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                                           // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                  // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                        // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                         // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                        // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                      // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                       // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                      // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                   // versionRom_s1_translator:uav_waitrequest -> versionRom_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] versionrom_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                    // versionRom_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> versionRom_s1_translator:uav_burstcount
	wire   [31:0] versionrom_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                     // versionRom_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> versionRom_s1_translator:uav_writedata
	wire   [17:0] versionrom_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                       // versionRom_s1_translator_avalon_universal_slave_0_agent:m0_address -> versionRom_s1_translator:uav_address
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                         // versionRom_s1_translator_avalon_universal_slave_0_agent:m0_write -> versionRom_s1_translator:uav_write
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                          // versionRom_s1_translator_avalon_universal_slave_0_agent:m0_lock -> versionRom_s1_translator:uav_lock
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                          // versionRom_s1_translator_avalon_universal_slave_0_agent:m0_read -> versionRom_s1_translator:uav_read
	wire   [31:0] versionrom_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                      // versionRom_s1_translator:uav_readdata -> versionRom_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                 // versionRom_s1_translator:uav_readdatavalid -> versionRom_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                   // versionRom_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> versionRom_s1_translator:uav_debugaccess
	wire    [3:0] versionrom_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                    // versionRom_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> versionRom_s1_translator:uav_byteenable
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                            // versionRom_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                  // versionRom_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                          // versionRom_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                   // versionRom_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                  // versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> versionRom_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                         // versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> versionRom_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                               // versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> versionRom_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                       // versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> versionRom_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                // versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> versionRom_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                               // versionRom_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                             // versionRom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> versionRom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] versionrom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                              // versionRom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> versionRom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                             // versionRom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> versionRom_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cheri_avalon_master_0_translator_avalon_universal_master_0_waitrequest;                                                   // CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_waitrequest -> CHERI_avalon_master_0_translator:uav_waitrequest
	wire    [5:0] cheri_avalon_master_0_translator_avalon_universal_master_0_burstcount;                                                    // CHERI_avalon_master_0_translator:uav_burstcount -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [255:0] cheri_avalon_master_0_translator_avalon_universal_master_0_writedata;                                                     // CHERI_avalon_master_0_translator:uav_writedata -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cheri_avalon_master_0_translator_avalon_universal_master_0_address;                                                       // CHERI_avalon_master_0_translator:uav_address -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_address
	wire          cheri_avalon_master_0_translator_avalon_universal_master_0_lock;                                                          // CHERI_avalon_master_0_translator:uav_lock -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_lock
	wire          cheri_avalon_master_0_translator_avalon_universal_master_0_write;                                                         // CHERI_avalon_master_0_translator:uav_write -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_write
	wire          cheri_avalon_master_0_translator_avalon_universal_master_0_read;                                                          // CHERI_avalon_master_0_translator:uav_read -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_read
	wire  [255:0] cheri_avalon_master_0_translator_avalon_universal_master_0_readdata;                                                      // CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_readdata -> CHERI_avalon_master_0_translator:uav_readdata
	wire          cheri_avalon_master_0_translator_avalon_universal_master_0_debugaccess;                                                   // CHERI_avalon_master_0_translator:uav_debugaccess -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [31:0] cheri_avalon_master_0_translator_avalon_universal_master_0_byteenable;                                                    // CHERI_avalon_master_0_translator:uav_byteenable -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cheri_avalon_master_0_translator_avalon_universal_master_0_readdatavalid;                                                 // CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:av_readdatavalid -> CHERI_avalon_master_0_translator:uav_readdatavalid
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                            // peripheral_bridge_s0_translator:uav_waitrequest -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                             // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> peripheral_bridge_s0_translator:uav_burstcount
	wire   [31:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                              // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> peripheral_bridge_s0_translator:uav_writedata
	wire   [31:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                                                // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> peripheral_bridge_s0_translator:uav_address
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                                                  // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> peripheral_bridge_s0_translator:uav_write
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                                   // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> peripheral_bridge_s0_translator:uav_lock
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                                                   // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> peripheral_bridge_s0_translator:uav_read
	wire   [31:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                               // peripheral_bridge_s0_translator:uav_readdata -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                          // peripheral_bridge_s0_translator:uav_readdatavalid -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                            // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> peripheral_bridge_s0_translator:uav_debugaccess
	wire    [3:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                             // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> peripheral_bridge_s0_translator:uav_byteenable
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                     // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                                           // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                   // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                                            // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                                           // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                  // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                        // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                         // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                        // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                      // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                       // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                      // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                                           // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                                                 // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                                         // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [100:0] peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                                                  // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                                                 // addr_router:sink_ready -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                         // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [100:0] mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_data;                                          // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router:sink_ready -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                          // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [100:0] mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_data;                                           // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_001:sink_ready -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                           // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                 // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                         // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [100:0] onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                  // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                 // id_router_002:sink_ready -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                                  // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_valid;                                        // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                                // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire   [90:0] mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_data;                                         // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_ready;                                        // addr_router_001:sink_ready -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                   // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire   [90:0] altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                    // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                         // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                               // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                       // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire   [90:0] leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                               // id_router_004:sink_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                     // Switches_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                           // Switches_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                   // Switches_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire   [90:0] switches_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                            // Switches_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                           // id_router_005:sink_ready -> Switches_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [90:0] transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_data;                                                       // transmit_fifo_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_006:sink_ready -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                            // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                                  // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                          // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [90:0] transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                                   // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                                  // id_router_007:sink_ready -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // receive_fifo_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // receive_fifo_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // receive_fifo_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [90:0] receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_data;                                                       // receive_fifo_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_008:sink_ready -> receive_fifo_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                            // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                                  // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                          // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire   [90:0] receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_data;                                                   // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                                  // id_router_009:sink_ready -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                   // versionRom_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                         // versionRom_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                 // versionRom_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire   [90:0] versionrom_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                          // versionRom_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          versionrom_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                         // id_router_010:sink_ready -> versionRom_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_endofpacket;                                          // CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_valid;                                                // CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_startofpacket;                                        // CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [358:0] cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_data;                                                 // CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_ready;                                                // addr_router_002:sink_ready -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:cp_ready
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                            // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                                  // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                          // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [106:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                                                   // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                                  // id_router_011:sink_ready -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                                              // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                                    // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                                            // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [100:0] addr_router_src_data;                                                                                                     // addr_router:src_data -> limiter:cmd_sink_data
	wire    [2:0] addr_router_src_channel;                                                                                                  // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                                    // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                                              // limiter:rsp_src_endofpacket -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                                    // limiter:rsp_src_valid -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                                            // limiter:rsp_src_startofpacket -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [100:0] limiter_rsp_src_data;                                                                                                     // limiter:rsp_src_data -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [2:0] limiter_rsp_src_channel;                                                                                                  // limiter:rsp_src_channel -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                                    // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                                          // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                                // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                                        // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire   [90:0] addr_router_001_src_data;                                                                                                 // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire    [7:0] addr_router_001_src_channel;                                                                                              // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                                                // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                                          // limiter_001:rsp_src_endofpacket -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                                                // limiter_001:rsp_src_valid -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                                        // limiter_001:rsp_src_startofpacket -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [90:0] limiter_001_rsp_src_data;                                                                                                 // limiter_001:rsp_src_data -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [7:0] limiter_001_rsp_src_channel;                                                                                              // limiter_001:rsp_src_channel -> mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                                                // mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                                        // burst_adapter:source0_endofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                              // burst_adapter:source0_valid -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                                      // burst_adapter:source0_startofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] burst_adapter_source0_data;                                                                                               // burst_adapter:source0_data -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                              // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire          burst_adapter_source0_channel;                                                                                            // burst_adapter:source0_channel -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                           // rst_controller:reset_out -> [CHERI:csi_clockreset_reset_n, CHERI_avalon_master_0_translator:reset, CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:reset, addr_router:reset, addr_router_002:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_002:reset, dc_fifo_0:in_reset_n, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_011:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, limiter:reset, limiter_pipeline:reset, limiter_pipeline_001:reset, mkMTL_Framebuffer_Flash_0:csi_clockreset_reset_n, mkMTL_Framebuffer_Flash_0_s0_translator:reset, mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:reset, mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mm_clock_crossing_bridge_0:s0_reset, mm_clock_crossing_bridge_0_s0_translator:reset, mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:reset, mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory_MIPS:reset, onchip_memory_MIPS_s1_translator:reset, onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, peripheral_bridge:reset, peripheral_bridge_m0_translator:reset, peripheral_bridge_m0_translator_avalon_universal_master_0_agent:reset, peripheral_bridge_s0_translator:reset, peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:reset, peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_011:reset, rsp_xbar_mux:reset, width_adapter:reset, width_adapter_001:reset]
	wire          rst_controller_001_reset_out_reset;                                                                                       // rst_controller_001:reset_out -> [Altera_UP_SD_Card_Avalon_Interface_1:i_reset_n, Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator:reset, Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, AvalonStream2MTL_LCD24bit_0:csi_clockreset_reset_n, LEDs:reset_n, LEDs_s1_translator:reset, LEDs_s1_translator_avalon_universal_slave_0_agent:reset, LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Switches:reset_n, Switches_s1_translator:reset, Switches_s1_translator_avalon_universal_slave_0_agent:reset, Switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router_001:reset, cmd_xbar_demux_001:reset, dc_fifo_0:out_reset_n, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, limiter_001:reset, limiter_pipeline_002:reset, limiter_pipeline_003:reset, mm_clock_crossing_bridge_0:m0_reset, mm_clock_crossing_bridge_0_m0_translator:reset, mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent:reset, receive_fifo:rdreset_n, receive_fifo:wrreset_n, receive_fifo_out_csr_translator:reset, receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:reset, receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, receive_fifo_out_translator:reset, receive_fifo_out_translator_avalon_universal_slave_0_agent:reset, receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_mux_001:reset, timing_adapter:reset_n, timing_adapter_1:reset_n, transmit_fifo:reset_n, transmit_fifo_in_csr_translator:reset, transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:reset, transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, transmit_fifo_in_translator:reset, transmit_fifo_in_translator_avalon_universal_slave_0_agent:reset, transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, versionRom:reset, versionRom_s1_translator:reset, versionRom_s1_translator_avalon_universal_slave_0_agent:reset, versionRom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                          // cmd_xbar_demux:src0_endofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                                // cmd_xbar_demux:src0_valid -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                                        // cmd_xbar_demux:src0_startofpacket -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_src0_data;                                                                                                 // cmd_xbar_demux:src0_data -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_src0_channel;                                                                                              // cmd_xbar_demux:src0_channel -> mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                          // cmd_xbar_demux:src1_endofpacket -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                                // cmd_xbar_demux:src1_valid -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                                        // cmd_xbar_demux:src1_startofpacket -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_src1_data;                                                                                                 // cmd_xbar_demux:src1_data -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_src1_channel;                                                                                              // cmd_xbar_demux:src1_channel -> mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src2_endofpacket;                                                                                          // cmd_xbar_demux:src2_endofpacket -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                                // cmd_xbar_demux:src2_valid -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                                        // cmd_xbar_demux:src2_startofpacket -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_src2_data;                                                                                                 // cmd_xbar_demux:src2_data -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_src2_channel;                                                                                              // cmd_xbar_demux:src2_channel -> onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                          // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                                // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                                        // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [100:0] rsp_xbar_demux_src0_data;                                                                                                 // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [2:0] rsp_xbar_demux_src0_channel;                                                                                              // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                                // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                                      // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                            // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                                    // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [100:0] rsp_xbar_demux_001_src0_data;                                                                                             // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [2:0] rsp_xbar_demux_001_src0_channel;                                                                                          // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                            // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                                      // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                            // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                                    // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [100:0] rsp_xbar_demux_002_src0_data;                                                                                             // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [2:0] rsp_xbar_demux_002_src0_channel;                                                                                          // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                            // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_src0_ready;                                                                                                // mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire          id_router_src_endofpacket;                                                                                                // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                                      // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                              // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [100:0] id_router_src_data;                                                                                                       // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [2:0] id_router_src_channel;                                                                                                    // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                                      // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_demux_src1_ready;                                                                                                // mkMTL_Framebuffer_Flash_0_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire          id_router_001_src_endofpacket;                                                                                            // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                                  // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                          // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [100:0] id_router_001_src_data;                                                                                                   // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [2:0] id_router_001_src_channel;                                                                                                // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                                  // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_src2_ready;                                                                                                // onchip_memory_MIPS_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire          id_router_002_src_endofpacket;                                                                                            // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                                  // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                                          // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [100:0] id_router_002_src_data;                                                                                                   // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [2:0] id_router_002_src_channel;                                                                                                // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                                  // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                                      // cmd_xbar_demux_001:src0_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                            // cmd_xbar_demux_001:src0_valid -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                                    // cmd_xbar_demux_001:src0_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] cmd_xbar_demux_001_src0_data;                                                                                             // cmd_xbar_demux_001:src0_data -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_001_src0_channel;                                                                                          // cmd_xbar_demux_001:src0_channel -> Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                                      // cmd_xbar_demux_001:src1_endofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                            // cmd_xbar_demux_001:src1_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                                    // cmd_xbar_demux_001:src1_startofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] cmd_xbar_demux_001_src1_data;                                                                                             // cmd_xbar_demux_001:src1_data -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_001_src1_channel;                                                                                          // cmd_xbar_demux_001:src1_channel -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                                      // cmd_xbar_demux_001:src2_endofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                            // cmd_xbar_demux_001:src2_valid -> Switches_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                                    // cmd_xbar_demux_001:src2_startofpacket -> Switches_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] cmd_xbar_demux_001_src2_data;                                                                                             // cmd_xbar_demux_001:src2_data -> Switches_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_001_src2_channel;                                                                                          // cmd_xbar_demux_001:src2_channel -> Switches_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                                      // cmd_xbar_demux_001:src3_endofpacket -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                            // cmd_xbar_demux_001:src3_valid -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                                    // cmd_xbar_demux_001:src3_startofpacket -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] cmd_xbar_demux_001_src3_data;                                                                                             // cmd_xbar_demux_001:src3_data -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_001_src3_channel;                                                                                          // cmd_xbar_demux_001:src3_channel -> transmit_fifo_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                                      // cmd_xbar_demux_001:src4_endofpacket -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                            // cmd_xbar_demux_001:src4_valid -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                                    // cmd_xbar_demux_001:src4_startofpacket -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] cmd_xbar_demux_001_src4_data;                                                                                             // cmd_xbar_demux_001:src4_data -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_001_src4_channel;                                                                                          // cmd_xbar_demux_001:src4_channel -> transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                                      // cmd_xbar_demux_001:src5_endofpacket -> receive_fifo_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                                            // cmd_xbar_demux_001:src5_valid -> receive_fifo_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                                    // cmd_xbar_demux_001:src5_startofpacket -> receive_fifo_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] cmd_xbar_demux_001_src5_data;                                                                                             // cmd_xbar_demux_001:src5_data -> receive_fifo_out_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_001_src5_channel;                                                                                          // cmd_xbar_demux_001:src5_channel -> receive_fifo_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                                      // cmd_xbar_demux_001:src6_endofpacket -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                                            // cmd_xbar_demux_001:src6_valid -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                                    // cmd_xbar_demux_001:src6_startofpacket -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] cmd_xbar_demux_001_src6_data;                                                                                             // cmd_xbar_demux_001:src6_data -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_001_src6_channel;                                                                                          // cmd_xbar_demux_001:src6_channel -> receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                                      // cmd_xbar_demux_001:src7_endofpacket -> versionRom_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                                            // cmd_xbar_demux_001:src7_valid -> versionRom_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                                    // cmd_xbar_demux_001:src7_startofpacket -> versionRom_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] cmd_xbar_demux_001_src7_data;                                                                                             // cmd_xbar_demux_001:src7_data -> versionRom_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_001_src7_channel;                                                                                          // cmd_xbar_demux_001:src7_channel -> versionRom_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                                      // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                            // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                                    // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire   [90:0] rsp_xbar_demux_003_src0_data;                                                                                             // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink0_data
	wire    [7:0] rsp_xbar_demux_003_src0_channel;                                                                                          // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                            // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                                      // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                            // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                                    // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire   [90:0] rsp_xbar_demux_004_src0_data;                                                                                             // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink1_data
	wire    [7:0] rsp_xbar_demux_004_src0_channel;                                                                                          // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                            // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                                      // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                            // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                                    // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire   [90:0] rsp_xbar_demux_005_src0_data;                                                                                             // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink2_data
	wire    [7:0] rsp_xbar_demux_005_src0_channel;                                                                                          // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                            // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                                      // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                            // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                                    // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire   [90:0] rsp_xbar_demux_006_src0_data;                                                                                             // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink3_data
	wire    [7:0] rsp_xbar_demux_006_src0_channel;                                                                                          // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                            // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                                      // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                            // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                                    // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire   [90:0] rsp_xbar_demux_007_src0_data;                                                                                             // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink4_data
	wire    [7:0] rsp_xbar_demux_007_src0_channel;                                                                                          // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                            // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                                      // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                            // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                                    // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire   [90:0] rsp_xbar_demux_008_src0_data;                                                                                             // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink5_data
	wire    [7:0] rsp_xbar_demux_008_src0_channel;                                                                                          // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                            // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                                      // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                            // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                                    // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire   [90:0] rsp_xbar_demux_009_src0_data;                                                                                             // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink6_data
	wire    [7:0] rsp_xbar_demux_009_src0_channel;                                                                                          // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                            // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                                      // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                            // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                                    // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire   [90:0] rsp_xbar_demux_010_src0_data;                                                                                             // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink7_data
	wire    [7:0] rsp_xbar_demux_010_src0_channel;                                                                                          // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                            // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_010:src0_ready
	wire          cmd_xbar_demux_001_src0_ready;                                                                                            // Altera_UP_SD_Card_Avalon_Interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src0_ready
	wire          id_router_003_src_endofpacket;                                                                                            // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                                  // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                          // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire   [90:0] id_router_003_src_data;                                                                                                   // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [7:0] id_router_003_src_channel;                                                                                                // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                                  // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src1_ready;                                                                                            // LEDs_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src1_ready
	wire          id_router_004_src_endofpacket;                                                                                            // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                                  // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                          // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire   [90:0] id_router_004_src_data;                                                                                                   // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [7:0] id_router_004_src_channel;                                                                                                // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                                  // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src2_ready;                                                                                            // Switches_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire          id_router_005_src_endofpacket;                                                                                            // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                                  // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                                          // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire   [90:0] id_router_005_src_data;                                                                                                   // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire    [7:0] id_router_005_src_channel;                                                                                                // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                                  // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                                            // transmit_fifo_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_006_src_endofpacket;                                                                                            // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                                  // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                          // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [90:0] id_router_006_src_data;                                                                                                   // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire    [7:0] id_router_006_src_channel;                                                                                                // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                                  // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                                            // transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_007_src_endofpacket;                                                                                            // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                                  // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                          // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [90:0] id_router_007_src_data;                                                                                                   // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire    [7:0] id_router_007_src_channel;                                                                                                // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                                  // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                                            // receive_fifo_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_008_src_endofpacket;                                                                                            // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                                  // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                          // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [90:0] id_router_008_src_data;                                                                                                   // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire    [7:0] id_router_008_src_channel;                                                                                                // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                                  // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                                            // receive_fifo_out_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_009_src_endofpacket;                                                                                            // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                                  // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                          // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire   [90:0] id_router_009_src_data;                                                                                                   // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire    [7:0] id_router_009_src_channel;                                                                                                // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                                  // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                                            // versionRom_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_010_src_endofpacket;                                                                                            // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                                  // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                                          // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire   [90:0] id_router_010_src_data;                                                                                                   // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire    [7:0] id_router_010_src_channel;                                                                                                // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                                  // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                                      // cmd_xbar_demux_002:src0_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                                            // cmd_xbar_demux_002:src0_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                                    // cmd_xbar_demux_002:src0_startofpacket -> width_adapter:in_startofpacket
	wire  [358:0] cmd_xbar_demux_002_src0_data;                                                                                             // cmd_xbar_demux_002:src0_data -> width_adapter:in_data
	wire    [0:0] cmd_xbar_demux_002_src0_channel;                                                                                          // cmd_xbar_demux_002:src0_channel -> width_adapter:in_channel
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                                      // rsp_xbar_demux_011:src0_endofpacket -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                            // rsp_xbar_demux_011:src0_valid -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                                    // rsp_xbar_demux_011:src0_startofpacket -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [358:0] rsp_xbar_demux_011_src0_data;                                                                                             // rsp_xbar_demux_011:src0_data -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:rp_data
	wire    [0:0] rsp_xbar_demux_011_src0_channel;                                                                                          // rsp_xbar_demux_011:src0_channel -> CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_002_src_endofpacket;                                                                                          // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                                // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                                        // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [358:0] addr_router_002_src_data;                                                                                                 // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [0:0] addr_router_002_src_channel;                                                                                              // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                                // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_011_src0_ready;                                                                                            // CHERI_avalon_master_0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_011:src0_ready
	wire          cmd_xbar_demux_002_src0_ready;                                                                                            // width_adapter:in_ready -> cmd_xbar_demux_002:src0_ready
	wire          width_adapter_src_endofpacket;                                                                                            // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                                  // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                                          // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [106:0] width_adapter_src_data;                                                                                                   // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                                                  // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire          width_adapter_src_channel;                                                                                                // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_011_src_endofpacket;                                                                                            // id_router_011:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_011_src_valid;                                                                                                  // id_router_011:src_valid -> width_adapter_001:in_valid
	wire          id_router_011_src_startofpacket;                                                                                          // id_router_011:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [106:0] id_router_011_src_data;                                                                                                   // id_router_011:src_data -> width_adapter_001:in_data
	wire    [0:0] id_router_011_src_channel;                                                                                                // id_router_011:src_channel -> width_adapter_001:in_channel
	wire          id_router_011_src_ready;                                                                                                  // width_adapter_001:in_ready -> id_router_011:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                                        // width_adapter_001:out_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                                              // width_adapter_001:out_valid -> rsp_xbar_demux_011:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                                      // width_adapter_001:out_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [358:0] width_adapter_001_src_data;                                                                                               // width_adapter_001:out_data -> rsp_xbar_demux_011:sink_data
	wire          width_adapter_001_src_ready;                                                                                              // rsp_xbar_demux_011:sink_ready -> width_adapter_001:out_ready
	wire          width_adapter_001_src_channel;                                                                                            // width_adapter_001:out_channel -> rsp_xbar_demux_011:sink_channel
	wire          limiter_pipeline_source0_endofpacket;                                                                                     // limiter_pipeline:out_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_pipeline_source0_valid;                                                                                           // limiter_pipeline:out_valid -> cmd_xbar_demux:sink_valid
	wire          limiter_pipeline_source0_startofpacket;                                                                                   // limiter_pipeline:out_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [100:0] limiter_pipeline_source0_data;                                                                                            // limiter_pipeline:out_data -> cmd_xbar_demux:sink_data
	wire    [2:0] limiter_pipeline_source0_channel;                                                                                         // limiter_pipeline:out_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_pipeline_source0_ready;                                                                                           // cmd_xbar_demux:sink_ready -> limiter_pipeline:out_ready
	wire          limiter_cmd_src_endofpacket;                                                                                              // limiter:cmd_src_endofpacket -> limiter_pipeline:in_endofpacket
	wire    [0:0] limiter_cmd_src_valid;                                                                                                    // limiter:cmd_src_valid -> limiter_pipeline:in_valid
	wire          limiter_cmd_src_startofpacket;                                                                                            // limiter:cmd_src_startofpacket -> limiter_pipeline:in_startofpacket
	wire  [100:0] limiter_cmd_src_data;                                                                                                     // limiter:cmd_src_data -> limiter_pipeline:in_data
	wire    [2:0] limiter_cmd_src_channel;                                                                                                  // limiter:cmd_src_channel -> limiter_pipeline:in_channel
	wire          limiter_cmd_src_ready;                                                                                                    // limiter_pipeline:in_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                             // rsp_xbar_mux:src_endofpacket -> limiter_pipeline_001:in_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                                   // rsp_xbar_mux:src_valid -> limiter_pipeline_001:in_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                           // rsp_xbar_mux:src_startofpacket -> limiter_pipeline_001:in_startofpacket
	wire  [100:0] rsp_xbar_mux_src_data;                                                                                                    // rsp_xbar_mux:src_data -> limiter_pipeline_001:in_data
	wire    [2:0] rsp_xbar_mux_src_channel;                                                                                                 // rsp_xbar_mux:src_channel -> limiter_pipeline_001:in_channel
	wire          rsp_xbar_mux_src_ready;                                                                                                   // limiter_pipeline_001:in_ready -> rsp_xbar_mux:src_ready
	wire          limiter_pipeline_001_source0_endofpacket;                                                                                 // limiter_pipeline_001:out_endofpacket -> limiter:rsp_sink_endofpacket
	wire          limiter_pipeline_001_source0_valid;                                                                                       // limiter_pipeline_001:out_valid -> limiter:rsp_sink_valid
	wire          limiter_pipeline_001_source0_startofpacket;                                                                               // limiter_pipeline_001:out_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [100:0] limiter_pipeline_001_source0_data;                                                                                        // limiter_pipeline_001:out_data -> limiter:rsp_sink_data
	wire    [2:0] limiter_pipeline_001_source0_channel;                                                                                     // limiter_pipeline_001:out_channel -> limiter:rsp_sink_channel
	wire          limiter_pipeline_001_source0_ready;                                                                                       // limiter:rsp_sink_ready -> limiter_pipeline_001:out_ready
	wire          limiter_pipeline_002_source0_endofpacket;                                                                                 // limiter_pipeline_002:out_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_pipeline_002_source0_valid;                                                                                       // limiter_pipeline_002:out_valid -> cmd_xbar_demux_001:sink_valid
	wire          limiter_pipeline_002_source0_startofpacket;                                                                               // limiter_pipeline_002:out_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire   [90:0] limiter_pipeline_002_source0_data;                                                                                        // limiter_pipeline_002:out_data -> cmd_xbar_demux_001:sink_data
	wire    [7:0] limiter_pipeline_002_source0_channel;                                                                                     // limiter_pipeline_002:out_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_pipeline_002_source0_ready;                                                                                       // cmd_xbar_demux_001:sink_ready -> limiter_pipeline_002:out_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                                          // limiter_001:cmd_src_endofpacket -> limiter_pipeline_002:in_endofpacket
	wire    [0:0] limiter_001_cmd_src_valid;                                                                                                // limiter_001:cmd_src_valid -> limiter_pipeline_002:in_valid
	wire          limiter_001_cmd_src_startofpacket;                                                                                        // limiter_001:cmd_src_startofpacket -> limiter_pipeline_002:in_startofpacket
	wire   [90:0] limiter_001_cmd_src_data;                                                                                                 // limiter_001:cmd_src_data -> limiter_pipeline_002:in_data
	wire    [7:0] limiter_001_cmd_src_channel;                                                                                              // limiter_001:cmd_src_channel -> limiter_pipeline_002:in_channel
	wire          limiter_001_cmd_src_ready;                                                                                                // limiter_pipeline_002:in_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                                         // rsp_xbar_mux_001:src_endofpacket -> limiter_pipeline_003:in_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                               // rsp_xbar_mux_001:src_valid -> limiter_pipeline_003:in_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                                       // rsp_xbar_mux_001:src_startofpacket -> limiter_pipeline_003:in_startofpacket
	wire   [90:0] rsp_xbar_mux_001_src_data;                                                                                                // rsp_xbar_mux_001:src_data -> limiter_pipeline_003:in_data
	wire    [7:0] rsp_xbar_mux_001_src_channel;                                                                                             // rsp_xbar_mux_001:src_channel -> limiter_pipeline_003:in_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                               // limiter_pipeline_003:in_ready -> rsp_xbar_mux_001:src_ready
	wire          limiter_pipeline_003_source0_endofpacket;                                                                                 // limiter_pipeline_003:out_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          limiter_pipeline_003_source0_valid;                                                                                       // limiter_pipeline_003:out_valid -> limiter_001:rsp_sink_valid
	wire          limiter_pipeline_003_source0_startofpacket;                                                                               // limiter_pipeline_003:out_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire   [90:0] limiter_pipeline_003_source0_data;                                                                                        // limiter_pipeline_003:out_data -> limiter_001:rsp_sink_data
	wire    [7:0] limiter_pipeline_003_source0_channel;                                                                                     // limiter_pipeline_003:out_channel -> limiter_001:rsp_sink_channel
	wire          limiter_pipeline_003_source0_ready;                                                                                       // limiter_001:rsp_sink_ready -> limiter_pipeline_003:out_ready
	wire    [4:0] cheri_irq_irq;                                                                                                            // irq_mapper:sender_irq -> CHERI:avm_irq_irqs
	wire          irq_mapper_receiver0_irq;                                                                                                 // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                                            // receive_fifo:rdclk_control_slave_irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver1_irq;                                                                                                 // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                                                        // transmit_fifo:wrclk_control_slave_irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver2_irq;                                                                                                 // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                                                                                        // Altera_UP_SD_Card_Avalon_Interface_1:o_avalon_irq -> irq_synchronizer_002:receiver_irq

	DE4_SOPC_onchip_memory_MIPS onchip_memory_mips (
		.clk        (clk_50),                                                          //   clk1.clk
		.address    (onchip_memory_mips_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory_mips_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory_mips_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory_mips_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory_mips_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory_mips_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory_mips_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                                   // reset1.reset
	);

	DE4_SOPC_LEDs leds (
		.clk        (clk_50),                                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address    (leds_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~leds_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (leds_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (leds_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (leds_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (leds_external_connection_export)                    // external_connection.export
	);

	mkTopAvalonPhy cheri (
		.csi_clockreset_clk                 (clk_50),                              //              clockreset.clk
		.csi_clockreset_reset_n             (~rst_controller_reset_out_reset),     //        clockreset_reset.reset_n
		.avm_readdata                       (cheri_avalon_master_0_readdata),      //         avalon_master_0.readdata
		.avm_readdatavalid                  (cheri_avalon_master_0_readdatavalid), //                        .readdatavalid
		.avm_waitrequest                    (cheri_avalon_master_0_waitrequest),   //                        .waitrequest
		.avm_writedata                      (cheri_avalon_master_0_writedata),     //                        .writedata
		.avm_address                        (cheri_avalon_master_0_address),       //                        .address
		.avm_read                           (cheri_avalon_master_0_read),          //                        .read
		.avm_write                          (cheri_avalon_master_0_write),         //                        .write
		.avm_byteenable                     (cheri_avalon_master_0_byteenable),    //                        .byteenable
		.avm_irq_irqs                       (cheri_irq_irq),                       //                     irq.irq
		.debugStreamSink_stream_in_data     (),                                    //   avalon_streaming_sink.data
		.debugStreamSink_stream_in_valid    (),                                    //                        .valid
		.debugStreamSource_stream_out_data  (),                                    // avalon_streaming_source.data
		.debugStreamSource_stream_out_valid (),                                    //                        .valid
		.debugStreamSource_stream_out_ready ()                                     //                        .ready
	);

	DE4_SOPC_transmit_fifo transmit_fifo (
		.wrclock                          (clk_50),                                                        //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),                           // reset_in.reset_n
		.avalonmm_write_slave_writedata   (transmit_fifo_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (transmit_fifo_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_address     (transmit_fifo_in_translator_avalon_anti_slave_0_address),       //         .address
		.avalonmm_write_slave_waitrequest (transmit_fifo_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (transmit_fifo_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (transmit_fifo_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (transmit_fifo_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (transmit_fifo_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (transmit_fifo_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_synchronizer_001_receiver_irq),                             //   in_irq.irq
		.avalonst_source_valid            (transmit_fifo_out_valid),                                       //      out.valid
		.avalonst_source_data             (transmit_fifo_out_data),                                        //         .data
		.avalonst_source_error            (transmit_fifo_out_error),                                       //         .error
		.avalonst_source_startofpacket    (transmit_fifo_out_startofpacket),                               //         .startofpacket
		.avalonst_source_endofpacket      (transmit_fifo_out_endofpacket),                                 //         .endofpacket
		.avalonst_source_empty            (transmit_fifo_out_empty),                                       //         .empty
		.avalonst_source_ready            (transmit_fifo_out_ready)                                        //         .ready
	);

	DE4_SOPC_receive_fifo receive_fifo (
		.wrclock                         (clk_50),                                                        //    clk_in.clk
		.wrreset_n                       (~rst_controller_001_reset_out_reset),                           //  reset_in.reset_n
		.avalonst_sink_valid             (timing_adapter_1_out_valid),                                    //        in.valid
		.avalonst_sink_data              (timing_adapter_1_out_data),                                     //          .data
		.avalonst_sink_error             (timing_adapter_1_out_error),                                    //          .error
		.avalonst_sink_startofpacket     (timing_adapter_1_out_startofpacket),                            //          .startofpacket
		.avalonst_sink_endofpacket       (timing_adapter_1_out_endofpacket),                              //          .endofpacket
		.avalonst_sink_empty             (timing_adapter_1_out_empty),                                    //          .empty
		.avalonst_sink_ready             (timing_adapter_1_out_ready),                                    //          .ready
		.rdclock                         (clk_50),                                                        //   clk_out.clk
		.rdreset_n                       (~rst_controller_001_reset_out_reset),                           // reset_out.reset_n
		.avalonmm_read_slave_readdata    (receive_fifo_out_translator_avalon_anti_slave_0_readdata),      //       out.readdata
		.avalonmm_read_slave_read        (receive_fifo_out_translator_avalon_anti_slave_0_read),          //          .read
		.avalonmm_read_slave_address     (receive_fifo_out_translator_avalon_anti_slave_0_address),       //          .address
		.avalonmm_read_slave_waitrequest (receive_fifo_out_translator_avalon_anti_slave_0_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address     (receive_fifo_out_csr_translator_avalon_anti_slave_0_address),   //   out_csr.address
		.rdclk_control_slave_read        (receive_fifo_out_csr_translator_avalon_anti_slave_0_read),      //          .read
		.rdclk_control_slave_writedata   (receive_fifo_out_csr_translator_avalon_anti_slave_0_writedata), //          .writedata
		.rdclk_control_slave_write       (receive_fifo_out_csr_translator_avalon_anti_slave_0_write),     //          .write
		.rdclk_control_slave_readdata    (receive_fifo_out_csr_translator_avalon_anti_slave_0_readdata),  //          .readdata
		.rdclk_control_slave_irq         (irq_synchronizer_receiver_irq)                                  //   out_irq.irq
	);

	DE4_SOPC_timing_adapter timing_adapter (
		.clk               (clk_50),                              //   clk.clk
		.reset_n           (~rst_controller_001_reset_out_reset), // reset.reset_n
		.in_ready          (transmit_fifo_out_ready),             //    in.ready
		.in_valid          (transmit_fifo_out_valid),             //      .valid
		.in_data           (transmit_fifo_out_data),              //      .data
		.in_error          (transmit_fifo_out_error),             //      .error
		.in_startofpacket  (transmit_fifo_out_startofpacket),     //      .startofpacket
		.in_endofpacket    (transmit_fifo_out_endofpacket),       //      .endofpacket
		.in_empty          (transmit_fifo_out_empty),             //      .empty
		.out_ready         (),                                    //   out.ready
		.out_valid         (),                                    //      .valid
		.out_data          (),                                    //      .data
		.out_error         (),                                    //      .error
		.out_startofpacket (),                                    //      .startofpacket
		.out_endofpacket   (),                                    //      .endofpacket
		.out_empty         ()                                     //      .empty
	);

	DE4_SOPC_timing_adapter_1 timing_adapter_1 (
		.clk               (clk_50),                              //   clk.clk
		.reset_n           (~rst_controller_001_reset_out_reset), // reset.reset_n
		.in_ready          (),                                    //    in.ready
		.in_valid          (),                                    //      .valid
		.in_data           (),                                    //      .data
		.in_error          (),                                    //      .error
		.in_startofpacket  (),                                    //      .startofpacket
		.in_endofpacket    (),                                    //      .endofpacket
		.in_empty          (),                                    //      .empty
		.out_ready         (timing_adapter_1_out_ready),          //   out.ready
		.out_valid         (timing_adapter_1_out_valid),          //      .valid
		.out_data          (timing_adapter_1_out_data),           //      .data
		.out_error         (timing_adapter_1_out_error),          //      .error
		.out_startofpacket (timing_adapter_1_out_startofpacket),  //      .startofpacket
		.out_endofpacket   (timing_adapter_1_out_endofpacket),    //      .endofpacket
		.out_empty         (timing_adapter_1_out_empty)           //      .empty
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (30),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) peripheral_bridge (
		.clk              (clk_50),                                                            //   clk.clk
		.reset            (rst_controller_reset_out_reset),                                    // reset.reset
		.s0_waitrequest   (peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.s0_readdatavalid (peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.s0_writedata     (peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.s0_address       (peripheral_bridge_s0_translator_avalon_anti_slave_0_address),       //      .address
		.s0_write         (peripheral_bridge_s0_translator_avalon_anti_slave_0_write),         //      .write
		.s0_read          (peripheral_bridge_s0_translator_avalon_anti_slave_0_read),          //      .read
		.s0_byteenable    (peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.s0_debugaccess   (peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (peripheral_bridge_m0_waitrequest),                                  //    m0.waitrequest
		.m0_readdata      (peripheral_bridge_m0_readdata),                                     //      .readdata
		.m0_readdatavalid (peripheral_bridge_m0_readdatavalid),                                //      .readdatavalid
		.m0_burstcount    (peripheral_bridge_m0_burstcount),                                   //      .burstcount
		.m0_writedata     (peripheral_bridge_m0_writedata),                                    //      .writedata
		.m0_address       (peripheral_bridge_m0_address),                                      //      .address
		.m0_write         (peripheral_bridge_m0_write),                                        //      .write
		.m0_read          (peripheral_bridge_m0_read),                                         //      .read
		.m0_byteenable    (peripheral_bridge_m0_byteenable),                                   //      .byteenable
		.m0_debugaccess   (peripheral_bridge_m0_debugaccess)                                   //      .debugaccess
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (24),
		.FIFO_DEPTH         (32),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (2),
		.RD_SYNC_DEPTH      (2)
	) dc_fifo_0 (
		.in_clk            (clk_50),                                             //        in_clk.clk
		.in_reset_n        (~rst_controller_reset_out_reset),                    //  in_clk_reset.reset_n
		.out_clk           (clk_50),                                             //       out_clk.clk
		.out_reset_n       (~rst_controller_001_reset_out_reset),                // out_clk_reset.reset_n
		.in_data           (mkmtl_framebuffer_flash_0_stream_out_data),          //            in.data
		.in_valid          (mkmtl_framebuffer_flash_0_stream_out_valid),         //              .valid
		.in_ready          (mkmtl_framebuffer_flash_0_stream_out_ready),         //              .ready
		.in_startofpacket  (mkmtl_framebuffer_flash_0_stream_out_startofpacket), //              .startofpacket
		.in_endofpacket    (mkmtl_framebuffer_flash_0_stream_out_endofpacket),   //              .endofpacket
		.out_data          (dc_fifo_0_out_data),                                 //           out.data
		.out_valid         (dc_fifo_0_out_valid),                                //              .valid
		.out_ready         (dc_fifo_0_out_ready),                                //              .ready
		.out_startofpacket (dc_fifo_0_out_startofpacket),                        //              .startofpacket
		.out_endofpacket   (dc_fifo_0_out_endofpacket),                          //              .endofpacket
		.in_csr_address    (1'b0),                                               //   (terminated)
		.in_csr_read       (1'b0),                                               //   (terminated)
		.in_csr_write      (1'b0),                                               //   (terminated)
		.in_csr_readdata   (),                                                   //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000),               //   (terminated)
		.out_csr_address   (1'b0),                                               //   (terminated)
		.out_csr_read      (1'b0),                                               //   (terminated)
		.out_csr_write     (1'b0),                                               //   (terminated)
		.out_csr_readdata  (),                                                   //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000)                //   (terminated)
	);

	mkAvalonStream2MTL_LCD24bit avalonstream2mtl_lcd24bit_0 (
		.csi_clockreset_clk          (clk_50),                              //       clockreset.clk
		.csi_clockreset_reset_n      (~rst_controller_001_reset_out_reset), // clockreset_reset.reset_n
		.asi_stream_in_data          (dc_fifo_0_out_data),                  //        stream_in.data
		.asi_stream_in_valid         (dc_fifo_0_out_valid),                 //                 .valid
		.asi_stream_in_startofpacket (dc_fifo_0_out_startofpacket),         //                 .startofpacket
		.asi_stream_in_endofpacket   (dc_fifo_0_out_endofpacket),           //                 .endofpacket
		.asi_stream_in_ready         (dc_fifo_0_out_ready),                 //                 .ready
		.coe_tpadlcd_mtl_r           (mtl_lcd_r),                           //    conduit_end_0.export
		.coe_tpadlcd_mtl_g           (mtl_lcd_g),                           //                 .export
		.coe_tpadlcd_mtl_b           (mtl_lcd_b),                           //                 .export
		.coe_tpadlcd_mtl_hsd         (mtl_lcd_hsd),                         //                 .export
		.coe_tpadlcd_mtl_vsd         (mtl_lcd_vsd)                          //                 .export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (18),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_0 (
		.m0_clk           (clk_50),                                                                     //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                                         // m0_reset.reset
		.s0_clk           (clk_50),                                                                     //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                                             // s0_reset.reset
		.s0_waitrequest   (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_0_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_0_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_0_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_0_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_0_m0_writedata),                                    //         .writedata
		.m0_address       (mm_clock_crossing_bridge_0_m0_address),                                      //         .address
		.m0_write         (mm_clock_crossing_bridge_0_m0_write),                                        //         .write
		.m0_read          (mm_clock_crossing_bridge_0_m0_read),                                         //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_0_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_0_m0_debugaccess)                                   //         .debugaccess
	);

	mkMTL_Framebuffer_Flash mkmtl_framebuffer_flash_0 (
		.csi_clockreset_clk           (clk_50),                                                                  //        clockreset.clk
		.csi_clockreset_reset_n       (~rst_controller_reset_out_reset),                                         //  clockreset_reset.reset_n
		.avs_s0_address               (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_address),     //                s0.address
		.avs_s0_writedata             (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.avs_s0_write                 (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_write),       //                  .write
		.avs_s0_read                  (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_read),        //                  .read
		.avs_s0_byteenable            (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_byteenable),  //                  .byteenable
		.avs_s0_readdata              (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.avs_s0_waitrequest           (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.aso_stream_out_data          (mkmtl_framebuffer_flash_0_stream_out_data),                               //        stream_out.data
		.aso_stream_out_valid         (mkmtl_framebuffer_flash_0_stream_out_valid),                              //                  .valid
		.aso_stream_out_ready         (mkmtl_framebuffer_flash_0_stream_out_ready),                              //                  .ready
		.aso_stream_out_startofpacket (mkmtl_framebuffer_flash_0_stream_out_startofpacket),                      //                  .startofpacket
		.aso_stream_out_endofpacket   (mkmtl_framebuffer_flash_0_stream_out_endofpacket),                        //                  .endofpacket
		.coe_touch_x1                 (touch_x1),                                                                // conduit_end_touch.export
		.coe_touch_y1                 (touch_y1),                                                                //                  .export
		.coe_touch_x2                 (touch_x2),                                                                //                  .export
		.coe_touch_y2                 (touch_y2),                                                                //                  .export
		.coe_touch_count_gesture      (touch_count_gesture),                                                     //                  .export
		.coe_touch_touch_valid        (touch_touch_valid),                                                       //                  .export
		.coe_ssram_adv                (mem_ssram_adv),                                                           //   conduit_end_mem.export
		.coe_ssram_bwa_n              (mem_ssram_bwa_n),                                                         //                  .export
		.coe_ssram_bwb_n              (mem_ssram_bwb_n),                                                         //                  .export
		.coe_ssram_ce_n               (mem_ssram_ce_n),                                                          //                  .export
		.coe_ssram_cke_n              (mem_ssram_cke_n),                                                         //                  .export
		.coe_ssram_oe_n               (mem_ssram_oe_n),                                                          //                  .export
		.coe_ssram_we_n               (mem_ssram_we_n),                                                          //                  .export
		.coe_fsm_a                    (mem_fsm_a),                                                               //                  .export
		.coe_fsm_d_out                (mem_fsm_d_out),                                                           //                  .export
		.coe_fsm_d_in                 (mem_fsm_d_in),                                                            //                  .export
		.coe_fsm_dout_req             (mem_fsm_dout_req),                                                        //                  .export
		.coe_flash_adv_n              (mem_flash_adv_n),                                                         //                  .export
		.coe_flash_ce_n               (mem_flash_ce_n),                                                          //                  .export
		.coe_flash_clk                (mem_flash_clk),                                                           //                  .export
		.coe_flash_oe_n               (mem_flash_oe_n),                                                          //                  .export
		.coe_flash_we_n               (mem_flash_we_n)                                                           //                  .export
	);

	Altera_UP_SD_Card_Avalon_Interface #(
		.ADDRESS_BUFFER   (8'b00000000),
		.ADDRESS_CID      (8'b10000000),
		.ADDRESS_CSD      (8'b10000100),
		.ADDRESS_OCR      (8'b10001000),
		.ADDRESS_SR       (8'b10001001),
		.ADDRESS_RCA      (8'b10001010),
		.ADDRESS_ARGUMENT (8'b10001011),
		.ADDRESS_COMMAND  (8'b10001100),
		.ADDRESS_ASR      (8'b10001101),
		.ADDRESS_R1       (8'b10001110)
	) altera_up_sd_card_avalon_interface_1 (
		.i_avalon_chip_select (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),  //   avalon_slave_0.chipselect
		.o_avalon_readdata    (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //                 .readdata
		.i_avalon_writedata   (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //                 .writedata
		.i_avalon_byteenable  (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),  //                 .byteenable
		.i_avalon_write       (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_write),       //                 .write
		.i_avalon_read        (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_read),        //                 .read
		.i_avalon_address     (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_address),     //                 .address
		.o_avalon_waitrequest (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest), //                 .waitrequest
		.b_SD_cmd             (sd_b_SD_cmd),                                                                                    //      conduit_end.export
		.b_SD_dat             (sd_b_SD_dat),                                                                                    //                 .export
		.b_SD_dat3            (sd_b_SD_dat3),                                                                                   //                 .export
		.o_SD_clock           (sd_o_SD_clock),                                                                                  //                 .export
		.i_clock              (clk_50),                                                                                         //       clock_sink.clk
		.o_avalon_irq         (irq_synchronizer_002_receiver_irq),                                                              // interrupt_sender.irq
		.i_reset_n            (~rst_controller_001_reset_out_reset)                                                             //       reset_sink.reset_n
	);

	DE4_SOPC_Switches switches (
		.clk      (clk_50),                                              //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address  (switches_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (switches_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (switches_export)                                      // external_connection.export
	);

	DE4_SOPC_versionRom versionrom (
		.clk         (clk_50),                                                   //   clk1.clk
		.address     (versionrom_s1_translator_avalon_anti_slave_0_address),     //     s1.address
		.chipselect  (versionrom_s1_translator_avalon_anti_slave_0_chipselect),  //       .chipselect
		.clken       (versionrom_s1_translator_avalon_anti_slave_0_clken),       //       .clken
		.readdata    (versionrom_s1_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.write       (versionrom_s1_translator_avalon_anti_slave_0_write),       //       .write
		.writedata   (versionrom_s1_translator_avalon_anti_slave_0_writedata),   //       .writedata
		.debugaccess (versionrom_s1_translator_avalon_anti_slave_0_debugaccess), //       .debugaccess
		.byteenable  (versionrom_s1_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.reset       (rst_controller_001_reset_out_reset)                        // reset1.reset
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (30),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (30),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) peripheral_bridge_m0_translator (
		.clk                   (clk_50),                                                                  //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                     reset.reset
		.uav_address           (peripheral_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (peripheral_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (peripheral_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (peripheral_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (peripheral_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (peripheral_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (peripheral_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (peripheral_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (peripheral_bridge_m0_read),                                               //                          .read
		.av_readdata           (peripheral_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (peripheral_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (peripheral_bridge_m0_write),                                              //                          .write
		.av_writedata          (peripheral_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (peripheral_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                    //               (terminated)
		.av_begintransfer      (1'b0),                                                                    //               (terminated)
		.av_chipselect         (1'b0),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                    //               (terminated)
		.uav_clken             (),                                                                        //               (terminated)
		.av_clken              (1'b1)                                                                     //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (30),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mm_clock_crossing_bridge_0_s0_translator (
		.clk                   (clk_50),                                                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (mm_clock_crossing_bridge_0_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_chipselect         (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (30),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mkmtl_framebuffer_flash_0_s0_translator (
		.clk                   (clk_50),                                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address           (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (mkmtl_framebuffer_flash_0_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_burstcount         (),                                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.av_chipselect         (),                                                                                        //              (terminated)
		.av_clken              (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_debugaccess        (),                                                                                        //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (30),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_mips_s1_translator (
		.clk                   (clk_50),                                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory_mips_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory_mips_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory_mips_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory_mips_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory_mips_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory_mips_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory_mips_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                 //              (terminated)
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (18),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (18),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) mm_clock_crossing_bridge_0_m0_translator (
		.clk                   (clk_50),                                                                           //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                               //                     reset.reset
		.uav_address           (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (mm_clock_crossing_bridge_0_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (mm_clock_crossing_bridge_0_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (mm_clock_crossing_bridge_0_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (mm_clock_crossing_bridge_0_m0_byteenable),                                         //                          .byteenable
		.av_read               (mm_clock_crossing_bridge_0_m0_read),                                               //                          .read
		.av_readdata           (mm_clock_crossing_bridge_0_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (mm_clock_crossing_bridge_0_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (mm_clock_crossing_bridge_0_m0_write),                                              //                          .write
		.av_writedata          (mm_clock_crossing_bridge_0_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (mm_clock_crossing_bridge_0_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                             //               (terminated)
		.av_begintransfer      (1'b0),                                                                             //               (terminated)
		.av_chipselect         (1'b0),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                             //               (terminated)
		.uav_clken             (),                                                                                 //               (terminated)
		.av_clken              (1'b1)                                                                              //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator (
		.clk                   (clk_50),                                                                                                         //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                                             //                    reset.reset
		.uav_address           (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                                                               //              (terminated)
		.av_burstcount         (),                                                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                                                               //              (terminated)
		.av_lock               (),                                                                                                               //              (terminated)
		.av_clken              (),                                                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                                                           //              (terminated)
		.av_debugaccess        (),                                                                                                               //              (terminated)
		.av_outputenable       ()                                                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leds_s1_translator (
		.clk                   (clk_50),                                                             //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address           (leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (leds_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (leds_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (leds_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switches_s1_translator (
		.clk                   (clk_50),                                                                 //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address           (switches_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (switches_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (switches_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (switches_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (switches_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (switches_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                       //              (terminated)
		.av_read               (),                                                                       //              (terminated)
		.av_writedata          (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_chipselect         (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) transmit_fifo_in_translator (
		.clk                   (clk_50),                                                                      //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address           (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (transmit_fifo_in_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (transmit_fifo_in_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_writedata          (transmit_fifo_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (transmit_fifo_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_read               (),                                                                            //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                        //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_chipselect         (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) transmit_fifo_in_csr_translator (
		.clk                   (clk_50),                                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                              //                    reset.reset
		.uav_address           (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (transmit_fifo_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (transmit_fifo_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (transmit_fifo_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (transmit_fifo_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (transmit_fifo_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) receive_fifo_out_translator (
		.clk                   (clk_50),                                                                      //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address           (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (receive_fifo_out_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_read               (receive_fifo_out_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (receive_fifo_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (receive_fifo_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_write              (),                                                                            //              (terminated)
		.av_writedata          (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_chipselect         (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) receive_fifo_out_csr_translator (
		.clk                   (clk_50),                                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                              //                    reset.reset
		.uav_address           (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (receive_fifo_out_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (receive_fifo_out_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (receive_fifo_out_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (receive_fifo_out_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (receive_fifo_out_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (18),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) versionrom_s1_translator (
		.clk                   (clk_50),                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address           (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (versionrom_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (versionrom_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (versionrom_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (versionrom_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (versionrom_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (versionrom_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (versionrom_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_debugaccess        (versionrom_s1_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (256),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (32),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (6),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (32),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cheri_avalon_master_0_translator (
		.clk                   (clk_50),                                                                   //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                     reset.reset
		.uav_address           (cheri_avalon_master_0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cheri_avalon_master_0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cheri_avalon_master_0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cheri_avalon_master_0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cheri_avalon_master_0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cheri_avalon_master_0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cheri_avalon_master_0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cheri_avalon_master_0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cheri_avalon_master_0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cheri_avalon_master_0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cheri_avalon_master_0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cheri_avalon_master_0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cheri_avalon_master_0_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cheri_avalon_master_0_byteenable),                                         //                          .byteenable
		.av_read               (cheri_avalon_master_0_read),                                               //                          .read
		.av_readdata           (cheri_avalon_master_0_readdata),                                           //                          .readdata
		.av_readdatavalid      (cheri_avalon_master_0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cheri_avalon_master_0_write),                                              //                          .write
		.av_writedata          (cheri_avalon_master_0_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                     //               (terminated)
		.av_begintransfer      (1'b0),                                                                     //               (terminated)
		.av_chipselect         (1'b0),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                     //               (terminated)
		.av_debugaccess        (1'b0),                                                                     //               (terminated)
		.uav_clken             (),                                                                         //               (terminated)
		.av_clken              (1'b1)                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (30),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) peripheral_bridge_s0_translator (
		.clk                   (clk_50),                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (peripheral_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (peripheral_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (peripheral_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_BEGIN_BURST           (85),
		.PKT_BURSTWRAP_H           (77),
		.PKT_BURSTWRAP_L           (75),
		.PKT_BURST_SIZE_H          (80),
		.PKT_BURST_SIZE_L          (78),
		.PKT_BURST_TYPE_H          (82),
		.PKT_BURST_TYPE_L          (81),
		.PKT_BYTE_CNT_H            (74),
		.PKT_BYTE_CNT_L            (72),
		.PKT_ADDR_H                (65),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (66),
		.PKT_TRANS_POSTED          (67),
		.PKT_TRANS_WRITE           (68),
		.PKT_TRANS_READ            (69),
		.PKT_TRANS_LOCK            (70),
		.PKT_TRANS_EXCLUSIVE       (71),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (89),
		.PKT_THREAD_ID_H           (91),
		.PKT_THREAD_ID_L           (91),
		.PKT_CACHE_H               (98),
		.PKT_CACHE_L               (95),
		.PKT_DATA_SIDEBAND_H       (84),
		.PKT_DATA_SIDEBAND_L       (84),
		.PKT_QOS_H                 (86),
		.PKT_QOS_L                 (86),
		.PKT_ADDR_SIDEBAND_H       (83),
		.PKT_ADDR_SIDEBAND_L       (83),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (3),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) peripheral_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (clk_50),                                                                           //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (peripheral_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (peripheral_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (peripheral_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (peripheral_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (85),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (65),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (66),
		.PKT_TRANS_POSTED          (67),
		.PKT_TRANS_WRITE           (68),
		.PKT_TRANS_READ            (69),
		.PKT_TRANS_LOCK            (70),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (77),
		.PKT_BURSTWRAP_L           (75),
		.PKT_BYTE_CNT_H            (74),
		.PKT_BYTE_CNT_L            (72),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (80),
		.PKT_BURST_SIZE_L          (78),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                                        //                .channel
		.rf_sink_ready           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (9),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (85),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (65),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (66),
		.PKT_TRANS_POSTED          (67),
		.PKT_TRANS_WRITE           (68),
		.PKT_TRANS_READ            (69),
		.PKT_TRANS_LOCK            (70),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (77),
		.PKT_BURSTWRAP_L           (75),
		.PKT_BYTE_CNT_H            (74),
		.PKT_BYTE_CNT_L            (72),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (80),
		.PKT_BURST_SIZE_L          (78),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                                       //                .channel
		.rf_sink_ready           (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (85),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (65),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (66),
		.PKT_TRANS_POSTED          (67),
		.PKT_TRANS_WRITE           (68),
		.PKT_TRANS_READ            (69),
		.PKT_TRANS_LOCK            (70),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (77),
		.PKT_BURSTWRAP_L           (75),
		.PKT_BYTE_CNT_H            (74),
		.PKT_BYTE_CNT_L            (72),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (80),
		.PKT_BURST_SIZE_L          (78),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                                //                .channel
		.rf_sink_ready           (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_BEGIN_BURST           (73),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.PKT_BURST_TYPE_H          (70),
		.PKT_BURST_TYPE_L          (69),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_TRANS_EXCLUSIVE       (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (81),
		.PKT_THREAD_ID_L           (81),
		.PKT_CACHE_H               (88),
		.PKT_CACHE_L               (85),
		.PKT_DATA_SIDEBAND_H       (72),
		.PKT_DATA_SIDEBAND_L       (72),
		.PKT_QOS_H                 (74),
		.PKT_QOS_L                 (74),
		.PKT_ADDR_SIDEBAND_H       (71),
		.PKT_ADDR_SIDEBAND_L       (71),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (8),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent (
		.clk              (clk_50),                                                                                    //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.av_address       (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                                 //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                                  //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                               //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                         //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                           //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                                  //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                                       //       clk_reset.reset
		.m0_address              (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src0_ready),                                                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src0_valid),                                                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src0_data),                                                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src0_startofpacket),                                                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src0_endofpacket),                                                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src0_channel),                                                                                          //                .channel
		.rf_sink_ready           (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                                       // clk_reset.reset
		.in_data           (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                                                     // (terminated)
		.csr_readdata      (),                                                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                     // (terminated)
		.almost_full_data  (),                                                                                                                         // (terminated)
		.almost_empty_data (),                                                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                                                     // (terminated)
		.out_empty         (),                                                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                                                     // (terminated)
		.out_error         (),                                                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                                                     // (terminated)
		.out_channel       ()                                                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src1_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src1_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src1_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src1_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src1_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src1_channel),                                              //                .channel
		.rf_sink_ready           (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) switches_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (switches_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switches_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switches_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switches_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switches_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                  //                .channel
		.rf_sink_ready           (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) transmit_fifo_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (transmit_fifo_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                       //                .channel
		.rf_sink_ready           (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                           //                .channel
		.rf_sink_ready           (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) receive_fifo_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (receive_fifo_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                       //                .channel
		.rf_sink_ready           (receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (receive_fifo_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (receive_fifo_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (receive_fifo_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (receive_fifo_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (receive_fifo_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (receive_fifo_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (receive_fifo_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (receive_fifo_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) receive_fifo_out_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                           //                .channel
		.rf_sink_ready           (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (73),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (53),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (54),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.PKT_TRANS_READ            (57),
		.PKT_TRANS_LOCK            (58),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (68),
		.PKT_BURST_SIZE_L          (66),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) versionrom_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (versionrom_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (versionrom_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (versionrom_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (versionrom_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (versionrom_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (versionrom_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                    //                .channel
		.rf_sink_ready           (versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (versionrom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (versionrom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (versionrom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (versionrom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (versionrom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (versionrom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (versionrom_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (versionrom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (352),
		.PKT_PROTECTION_L          (350),
		.PKT_BEGIN_BURST           (345),
		.PKT_BURSTWRAP_H           (337),
		.PKT_BURSTWRAP_L           (332),
		.PKT_BURST_SIZE_H          (340),
		.PKT_BURST_SIZE_L          (338),
		.PKT_BURST_TYPE_H          (342),
		.PKT_BURST_TYPE_L          (341),
		.PKT_BYTE_CNT_H            (331),
		.PKT_BYTE_CNT_L            (326),
		.PKT_ADDR_H                (319),
		.PKT_ADDR_L                (288),
		.PKT_TRANS_COMPRESSED_READ (320),
		.PKT_TRANS_POSTED          (321),
		.PKT_TRANS_WRITE           (322),
		.PKT_TRANS_READ            (323),
		.PKT_TRANS_LOCK            (324),
		.PKT_TRANS_EXCLUSIVE       (325),
		.PKT_DATA_H                (255),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (287),
		.PKT_BYTEEN_L              (256),
		.PKT_SRC_ID_H              (347),
		.PKT_SRC_ID_L              (347),
		.PKT_DEST_ID_H             (348),
		.PKT_DEST_ID_L             (348),
		.PKT_THREAD_ID_H           (349),
		.PKT_THREAD_ID_L           (349),
		.PKT_CACHE_H               (356),
		.PKT_CACHE_L               (353),
		.PKT_DATA_SIDEBAND_H       (344),
		.PKT_DATA_SIDEBAND_L       (344),
		.PKT_QOS_H                 (346),
		.PKT_QOS_L                 (346),
		.PKT_ADDR_SIDEBAND_H       (343),
		.PKT_ADDR_SIDEBAND_L       (343),
		.ST_DATA_W                 (359),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (6),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (63),
		.CACHE_VALUE               (4'b0000)
	) cheri_avalon_master_0_translator_avalon_universal_master_0_agent (
		.clk              (clk_50),                                                                            //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (cheri_avalon_master_0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cheri_avalon_master_0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cheri_avalon_master_0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cheri_avalon_master_0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cheri_avalon_master_0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cheri_avalon_master_0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cheri_avalon_master_0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cheri_avalon_master_0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cheri_avalon_master_0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cheri_avalon_master_0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cheri_avalon_master_0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_011_src0_valid),                                                     //        rp.valid
		.rp_data          (rsp_xbar_demux_011_src0_data),                                                      //          .data
		.rp_channel       (rsp_xbar_demux_011_src0_channel),                                                   //          .channel
		.rp_startofpacket (rsp_xbar_demux_011_src0_startofpacket),                                             //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),                                               //          .endofpacket
		.rp_ready         (rsp_xbar_demux_011_src0_ready)                                                      //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (95),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (96),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) peripheral_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                               //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                               //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                         //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                             //                .channel
		.rf_sink_ready           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (5),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	DE4_SOPC_addr_router addr_router (
		.sink_ready         (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_src_valid),                                                            //          .valid
		.src_data           (addr_router_src_data),                                                             //          .data
		.src_channel        (addr_router_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                       //          .endofpacket
	);

	DE4_SOPC_id_router id_router (
		.sink_ready         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mm_clock_crossing_bridge_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_src_valid),                                                                      //          .valid
		.src_data           (id_router_src_data),                                                                       //          .data
		.src_channel        (id_router_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                 //          .endofpacket
	);

	DE4_SOPC_id_router id_router_001 (
		.sink_ready         (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mkmtl_framebuffer_flash_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_001_src_valid),                                                                 //          .valid
		.src_data           (id_router_001_src_data),                                                                  //          .data
		.src_channel        (id_router_001_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                            //          .endofpacket
	);

	DE4_SOPC_id_router id_router_002 (
		.sink_ready         (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_mips_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                          //       src.ready
		.src_valid          (id_router_002_src_valid),                                                          //          .valid
		.src_data           (id_router_002_src_data),                                                           //          .data
		.src_channel        (id_router_002_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                     //          .endofpacket
	);

	DE4_SOPC_addr_router_001 addr_router_001 (
		.sink_ready         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mm_clock_crossing_bridge_0_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                                 //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                                 //          .valid
		.src_data           (addr_router_001_src_data),                                                                  //          .data
		.src_channel        (addr_router_001_src_channel),                                                               //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                            //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_003 (
		.sink_ready         (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altera_up_sd_card_avalon_interface_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                                             // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                                        //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                                        //          .valid
		.src_data           (id_router_003_src_data),                                                                                         //          .data
		.src_channel        (id_router_003_src_channel),                                                                                      //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                                                //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                                                   //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_004 (
		.sink_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                            //       src.ready
		.src_valid          (id_router_004_src_valid),                                            //          .valid
		.src_data           (id_router_004_src_data),                                             //          .data
		.src_channel        (id_router_004_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                       //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_005 (
		.sink_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switches_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                //       src.ready
		.src_valid          (id_router_005_src_valid),                                                //          .valid
		.src_data           (id_router_005_src_data),                                                 //          .data
		.src_channel        (id_router_005_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                           //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_006 (
		.sink_ready         (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (transmit_fifo_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                     //       src.ready
		.src_valid          (id_router_006_src_valid),                                                     //          .valid
		.src_data           (id_router_006_src_data),                                                      //          .data
		.src_channel        (id_router_006_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_007 (
		.sink_ready         (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (transmit_fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                         //       src.ready
		.src_valid          (id_router_007_src_valid),                                                         //          .valid
		.src_data           (id_router_007_src_data),                                                          //          .data
		.src_channel        (id_router_007_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                    //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_008 (
		.sink_ready         (receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (receive_fifo_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                     //       src.ready
		.src_valid          (id_router_008_src_valid),                                                     //          .valid
		.src_data           (id_router_008_src_data),                                                      //          .data
		.src_channel        (id_router_008_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_009 (
		.sink_ready         (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (receive_fifo_out_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                         //       src.ready
		.src_valid          (id_router_009_src_valid),                                                         //          .valid
		.src_data           (id_router_009_src_data),                                                          //          .data
		.src_channel        (id_router_009_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                    //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_010 (
		.sink_ready         (versionrom_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (versionrom_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (versionrom_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (versionrom_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (versionrom_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                  //       src.ready
		.src_valid          (id_router_010_src_valid),                                                  //          .valid
		.src_data           (id_router_010_src_data),                                                   //          .data
		.src_channel        (id_router_010_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                             //          .endofpacket
	);

	DE4_SOPC_addr_router_002 addr_router_002 (
		.sink_ready         (cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cheri_avalon_master_0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                         //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                         //          .valid
		.src_data           (addr_router_002_src_data),                                                          //          .data
		.src_channel        (addr_router_002_src_channel),                                                       //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                    //          .endofpacket
	);

	DE4_SOPC_id_router_011 id_router_011 (
		.sink_ready         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                         //       src.ready
		.src_valid          (id_router_011_src_valid),                                                         //          .valid
		.src_data           (id_router_011_src_data),                                                          //          .data
		.src_channel        (id_router_011_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                    //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (89),
		.PKT_TRANS_POSTED          (67),
		.PKT_TRANS_WRITE           (68),
		.MAX_OUTSTANDING_RESPONSES (12),
		.PIPELINED                 (0),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (3),
		.VALID_WIDTH               (1),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (74),
		.PKT_BYTE_CNT_L            (72),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_50),                                     //       clk.clk
		.reset                  (rst_controller_reset_out_reset),             // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),                      //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),                      //          .valid
		.cmd_sink_data          (addr_router_src_data),                       //          .data
		.cmd_sink_channel       (addr_router_src_channel),                    //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),              //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),                //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),                      //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),                       //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),                    //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),              //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),                //          .endofpacket
		.cmd_src_valid          (limiter_cmd_src_valid),                      //          .valid
		.rsp_sink_ready         (limiter_pipeline_001_source0_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (limiter_pipeline_001_source0_valid),         //          .valid
		.rsp_sink_channel       (limiter_pipeline_001_source0_channel),       //          .channel
		.rsp_sink_data          (limiter_pipeline_001_source0_data),          //          .data
		.rsp_sink_startofpacket (limiter_pipeline_001_source0_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (limiter_pipeline_001_source0_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),                      //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),                      //          .valid
		.rsp_src_data           (limiter_rsp_src_data),                       //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),                    //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),              //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket)                 //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (78),
		.PKT_TRANS_POSTED          (55),
		.PKT_TRANS_WRITE           (56),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (8),
		.VALID_WIDTH               (1),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_50),                                     //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset),         // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),                  //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),                  //          .valid
		.cmd_sink_data          (addr_router_001_src_data),                   //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),                //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),          //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),            //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),                  //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),                   //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),                //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),          //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),            //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_src_valid),                  //          .valid
		.rsp_sink_ready         (limiter_pipeline_003_source0_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (limiter_pipeline_003_source0_valid),         //          .valid
		.rsp_sink_channel       (limiter_pipeline_003_source0_channel),       //          .channel
		.rsp_sink_data          (limiter_pipeline_003_source0_data),          //          .data
		.rsp_sink_startofpacket (limiter_pipeline_003_source0_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (limiter_pipeline_003_source0_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),                  //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),                  //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),                   //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),                //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),          //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket)             //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (93),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (1),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (85),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (63),
		.BURSTWRAP_CONST_VALUE     (63)
	) burst_adapter (
		.clk                   (clk_50),                              //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_50),                         //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_50),                             //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	DE4_SOPC_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_50),                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready         (limiter_pipeline_source0_ready),         //      sink.ready
		.sink_channel       (limiter_pipeline_source0_channel),       //          .channel
		.sink_data          (limiter_pipeline_source0_data),          //          .data
		.sink_startofpacket (limiter_pipeline_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (limiter_pipeline_source0_endofpacket),   //          .endofpacket
		.sink_valid         (limiter_pipeline_source0_valid),         //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),              //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),              //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),               //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),            //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),        //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),              //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),              //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),               //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),            //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),      //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),        //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),              //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),              //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),               //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),            //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),      //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)         //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_50),                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_50),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_50),                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),         // clk_reset.reset
		.sink_ready         (limiter_pipeline_002_source0_ready),         //      sink.ready
		.sink_channel       (limiter_pipeline_002_source0_channel),       //          .channel
		.sink_data          (limiter_pipeline_002_source0_data),          //          .data
		.sink_startofpacket (limiter_pipeline_002_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (limiter_pipeline_002_source0_endofpacket),   //          .endofpacket
		.sink_valid         (limiter_pipeline_002_source0_valid),         //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),              //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),              //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),               //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),            //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),        //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),              //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),              //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),               //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),            //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket),      //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),        //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),              //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),              //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),               //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),            //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket),      //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),        //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),              //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),              //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),               //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),            //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket),      //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),        //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),              //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),              //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),               //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),            //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket),      //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),        //          .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),              //      src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),              //          .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),               //          .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),            //          .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket),      //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),        //          .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),              //      src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),              //          .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),               //          .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),            //          .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket),      //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),        //          .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),              //      src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),              //          .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),               //          .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),            //          .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket),      //          .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)         //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_003 rsp_xbar_demux_006 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_003 rsp_xbar_demux_007 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_003 rsp_xbar_demux_008 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_003 rsp_xbar_demux_009 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_003 rsp_xbar_demux_010 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_50),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_003_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_004_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_005_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_006_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_007_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_008_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_009_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_010_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_002 rsp_xbar_demux_011 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (319),
		.IN_PKT_ADDR_L                 (288),
		.IN_PKT_DATA_H                 (255),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (287),
		.IN_PKT_BYTEEN_L               (256),
		.IN_PKT_BYTE_CNT_H             (331),
		.IN_PKT_BYTE_CNT_L             (326),
		.IN_PKT_TRANS_COMPRESSED_READ  (320),
		.IN_PKT_BURSTWRAP_H            (337),
		.IN_PKT_BURSTWRAP_L            (332),
		.IN_PKT_BURST_SIZE_H           (340),
		.IN_PKT_BURST_SIZE_L           (338),
		.IN_PKT_RESPONSE_STATUS_H      (358),
		.IN_PKT_RESPONSE_STATUS_L      (357),
		.IN_PKT_TRANS_EXCLUSIVE        (325),
		.IN_PKT_BURST_TYPE_H           (342),
		.IN_PKT_BURST_TYPE_L           (341),
		.IN_ST_DATA_W                  (359),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (79),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (88),
		.OUT_PKT_BURST_SIZE_L          (86),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (90),
		.OUT_PKT_BURST_TYPE_L          (89),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (clk_50),                                //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_002_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),         //       src.endofpacket
		.out_data             (width_adapter_src_data),                //          .data
		.out_channel          (width_adapter_src_channel),             //          .channel
		.out_valid            (width_adapter_src_valid),               //          .valid
		.out_ready            (width_adapter_src_ready),               //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),       //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (79),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (85),
		.IN_PKT_BURSTWRAP_L            (80),
		.IN_PKT_BURST_SIZE_H           (88),
		.IN_PKT_BURST_SIZE_L           (86),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (90),
		.IN_PKT_BURST_TYPE_L           (89),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (319),
		.OUT_PKT_ADDR_L                (288),
		.OUT_PKT_DATA_H                (255),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (287),
		.OUT_PKT_BYTEEN_L              (256),
		.OUT_PKT_BYTE_CNT_H            (331),
		.OUT_PKT_BYTE_CNT_L            (326),
		.OUT_PKT_TRANS_COMPRESSED_READ (320),
		.OUT_PKT_BURST_SIZE_H          (340),
		.OUT_PKT_BURST_SIZE_L          (338),
		.OUT_PKT_RESPONSE_STATUS_H     (358),
		.OUT_PKT_RESPONSE_STATUS_L     (357),
		.OUT_PKT_TRANS_EXCLUSIVE       (325),
		.OUT_PKT_BURST_TYPE_H          (342),
		.OUT_PKT_BURST_TYPE_L          (341),
		.OUT_ST_DATA_W                 (359),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (clk_50),                              //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_011_src_valid),             //      sink.valid
		.in_channel           (id_router_011_src_channel),           //          .channel
		.in_startofpacket     (id_router_011_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_011_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_011_src_ready),             //          .ready
		.in_data              (id_router_011_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (101),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) limiter_pipeline (
		.clk               (clk_50),                                 //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (limiter_cmd_src_ready),                  //     sink0.ready
		.in_valid          (limiter_cmd_src_valid),                  //          .valid
		.in_startofpacket  (limiter_cmd_src_startofpacket),          //          .startofpacket
		.in_endofpacket    (limiter_cmd_src_endofpacket),            //          .endofpacket
		.in_data           (limiter_cmd_src_data),                   //          .data
		.in_channel        (limiter_cmd_src_channel),                //          .channel
		.out_ready         (limiter_pipeline_source0_ready),         //   source0.ready
		.out_valid         (limiter_pipeline_source0_valid),         //          .valid
		.out_startofpacket (limiter_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (limiter_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (limiter_pipeline_source0_data),          //          .data
		.out_channel       (limiter_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (101),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) limiter_pipeline_001 (
		.clk               (clk_50),                                     //       cr0.clk
		.reset             (rst_controller_reset_out_reset),             // cr0_reset.reset
		.in_ready          (rsp_xbar_mux_src_ready),                     //     sink0.ready
		.in_valid          (rsp_xbar_mux_src_valid),                     //          .valid
		.in_startofpacket  (rsp_xbar_mux_src_startofpacket),             //          .startofpacket
		.in_endofpacket    (rsp_xbar_mux_src_endofpacket),               //          .endofpacket
		.in_data           (rsp_xbar_mux_src_data),                      //          .data
		.in_channel        (rsp_xbar_mux_src_channel),                   //          .channel
		.out_ready         (limiter_pipeline_001_source0_ready),         //   source0.ready
		.out_valid         (limiter_pipeline_001_source0_valid),         //          .valid
		.out_startofpacket (limiter_pipeline_001_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (limiter_pipeline_001_source0_endofpacket),   //          .endofpacket
		.out_data          (limiter_pipeline_001_source0_data),          //          .data
		.out_channel       (limiter_pipeline_001_source0_channel),       //          .channel
		.in_empty          (1'b0),                                       // (terminated)
		.out_empty         (),                                           // (terminated)
		.out_error         (),                                           // (terminated)
		.in_error          (1'b0)                                        // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (91),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (8),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) limiter_pipeline_002 (
		.clk               (clk_50),                                     //       cr0.clk
		.reset             (rst_controller_001_reset_out_reset),         // cr0_reset.reset
		.in_ready          (limiter_001_cmd_src_ready),                  //     sink0.ready
		.in_valid          (limiter_001_cmd_src_valid),                  //          .valid
		.in_startofpacket  (limiter_001_cmd_src_startofpacket),          //          .startofpacket
		.in_endofpacket    (limiter_001_cmd_src_endofpacket),            //          .endofpacket
		.in_data           (limiter_001_cmd_src_data),                   //          .data
		.in_channel        (limiter_001_cmd_src_channel),                //          .channel
		.out_ready         (limiter_pipeline_002_source0_ready),         //   source0.ready
		.out_valid         (limiter_pipeline_002_source0_valid),         //          .valid
		.out_startofpacket (limiter_pipeline_002_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (limiter_pipeline_002_source0_endofpacket),   //          .endofpacket
		.out_data          (limiter_pipeline_002_source0_data),          //          .data
		.out_channel       (limiter_pipeline_002_source0_channel),       //          .channel
		.in_empty          (1'b0),                                       // (terminated)
		.out_empty         (),                                           // (terminated)
		.out_error         (),                                           // (terminated)
		.in_error          (1'b0)                                        // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (91),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (8),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) limiter_pipeline_003 (
		.clk               (clk_50),                                     //       cr0.clk
		.reset             (rst_controller_001_reset_out_reset),         // cr0_reset.reset
		.in_ready          (rsp_xbar_mux_001_src_ready),                 //     sink0.ready
		.in_valid          (rsp_xbar_mux_001_src_valid),                 //          .valid
		.in_startofpacket  (rsp_xbar_mux_001_src_startofpacket),         //          .startofpacket
		.in_endofpacket    (rsp_xbar_mux_001_src_endofpacket),           //          .endofpacket
		.in_data           (rsp_xbar_mux_001_src_data),                  //          .data
		.in_channel        (rsp_xbar_mux_001_src_channel),               //          .channel
		.out_ready         (limiter_pipeline_003_source0_ready),         //   source0.ready
		.out_valid         (limiter_pipeline_003_source0_valid),         //          .valid
		.out_startofpacket (limiter_pipeline_003_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (limiter_pipeline_003_source0_endofpacket),   //          .endofpacket
		.out_data          (limiter_pipeline_003_source0_data),          //          .data
		.out_channel       (limiter_pipeline_003_source0_channel),       //          .channel
		.in_empty          (1'b0),                                       // (terminated)
		.out_empty         (),                                           // (terminated)
		.out_error         (),                                           // (terminated)
		.in_error          (1'b0)                                        // (terminated)
	);

	DE4_SOPC_irq_mapper irq_mapper (
		.clk           (clk_50),                         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cheri_irq_irq)                   //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_50),                             //       receiver_clk.clk
		.sender_clk     (clk_50),                             //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_50),                             //       receiver_clk.clk
		.sender_clk     (clk_50),                             //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_50),                             //       receiver_clk.clk
		.sender_clk     (clk_50),                             //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	assign sram_clk_clk = clk_50;

endmodule
