module my_fir_h1_altr_st (clk, 
              rst, 
              data_in, 
              rdy_to_ld, 
              done, 
              fir_result); 
parameter DATA_WIDTH  = 16;
parameter COEF_WIDTH  = 9;
parameter ACCUM_WIDTH = 28;

input clk, rst;
input [DATA_WIDTH-1:0] data_in;
output rdy_to_ld;
wire rdy_to_ld;
wire rdy_int;
output done;
wire done;
wire done_int;
assign rdy_to_ld = 1'b1;
assign done = 1'b1;
output [ACCUM_WIDTH-1:0] fir_result;
wire addr_low;
assign addr_low = 1'b0;
wire clk_en;
assign clk_en = 1'b1;


//--- Parallel TDL Storage ---
wire inv_rst;
assign inv_rst = ~rst;
wire [15:0] tdl_0_n;
wire [15:0] tdl_1_n;
wire [15:0] tdl_2_n;
wire [15:0] tdl_3_n;
wire [15:0] tdl_4_n;
wire [15:0] tdl_5_n;
wire [15:0] tdl_6_n;


//--- TDL  ---
tdl_da_lc Utdldalc0n (.clk(clk), .clk_en(inv_rst), .data_in(data_in), .data_out(tdl_0_n) );
defparam Utdldalc0n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc1n (.clk(clk), .clk_en(clk_en), .data_in(tdl_0_n), .data_out(tdl_1_n) );
defparam Utdldalc1n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc2n (.clk(clk), .clk_en(clk_en), .data_in(tdl_1_n), .data_out(tdl_2_n) );
defparam Utdldalc2n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc3n (.clk(clk), .clk_en(clk_en), .data_in(tdl_2_n), .data_out(tdl_3_n) );
defparam Utdldalc3n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc4n (.clk(clk), .clk_en(clk_en), .data_in(tdl_3_n), .data_out(tdl_4_n) );
defparam Utdldalc4n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc5n (.clk(clk), .clk_en(clk_en), .data_in(tdl_4_n), .data_out(tdl_5_n) );
defparam Utdldalc5n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc6n (.clk(clk), .clk_en(clk_en), .data_in(tdl_5_n), .data_out(tdl_6_n) );
defparam Utdldalc6n.WIDTH = DATA_WIDTH;


// --- ROM LUTs ---- 
wire [8:0] lut_val_0_n_0_pp;
rom_lut Ur0_n_0_pp (.addr_in( {tdl_4_n[0],tdl_2_n[0],tdl_1_n[0],tdl_0_n[0] } ), .data_out( lut_val_0_n_0_pp[8:0]) ) ;
 defparam Ur0_n_0_pp.DATA_WIDTH = 9;
defparam Ur0_n_0_pp.C0 = 0;
defparam Ur0_n_0_pp.C1 = 497;
defparam Ur0_n_0_pp.C2 = 25;
defparam Ur0_n_0_pp.C3 = 10;
defparam Ur0_n_0_pp.C4 = 193;
defparam Ur0_n_0_pp.C5 = 178;
defparam Ur0_n_0_pp.C6 = 218;
defparam Ur0_n_0_pp.C7 = 203;
defparam Ur0_n_0_pp.C8 = 319;
defparam Ur0_n_0_pp.C9 = 304;
defparam Ur0_n_0_pp.CA = 344;
defparam Ur0_n_0_pp.CB = 329;
defparam Ur0_n_0_pp.CC = 0;
defparam Ur0_n_0_pp.CD = 497;
defparam Ur0_n_0_pp.CE = 25;
defparam Ur0_n_0_pp.CF = 10;
wire [8:0] lut_val_0_n_1_pp;
rom_lut Ur0_n_1_pp (.addr_in( {tdl_4_n[1],tdl_2_n[1],tdl_1_n[1],tdl_0_n[1] } ), .data_out( lut_val_0_n_1_pp[8:0]) ) ;
 defparam Ur0_n_1_pp.DATA_WIDTH = 9;
defparam Ur0_n_1_pp.C0 = 0;
defparam Ur0_n_1_pp.C1 = 497;
defparam Ur0_n_1_pp.C2 = 25;
defparam Ur0_n_1_pp.C3 = 10;
defparam Ur0_n_1_pp.C4 = 193;
defparam Ur0_n_1_pp.C5 = 178;
defparam Ur0_n_1_pp.C6 = 218;
defparam Ur0_n_1_pp.C7 = 203;
defparam Ur0_n_1_pp.C8 = 319;
defparam Ur0_n_1_pp.C9 = 304;
defparam Ur0_n_1_pp.CA = 344;
defparam Ur0_n_1_pp.CB = 329;
defparam Ur0_n_1_pp.CC = 0;
defparam Ur0_n_1_pp.CD = 497;
defparam Ur0_n_1_pp.CE = 25;
defparam Ur0_n_1_pp.CF = 10;
wire [8:0] lut_val_0_n_2_pp;
rom_lut Ur0_n_2_pp (.addr_in( {tdl_4_n[2],tdl_2_n[2],tdl_1_n[2],tdl_0_n[2] } ), .data_out( lut_val_0_n_2_pp[8:0]) ) ;
 defparam Ur0_n_2_pp.DATA_WIDTH = 9;
defparam Ur0_n_2_pp.C0 = 0;
defparam Ur0_n_2_pp.C1 = 497;
defparam Ur0_n_2_pp.C2 = 25;
defparam Ur0_n_2_pp.C3 = 10;
defparam Ur0_n_2_pp.C4 = 193;
defparam Ur0_n_2_pp.C5 = 178;
defparam Ur0_n_2_pp.C6 = 218;
defparam Ur0_n_2_pp.C7 = 203;
defparam Ur0_n_2_pp.C8 = 319;
defparam Ur0_n_2_pp.C9 = 304;
defparam Ur0_n_2_pp.CA = 344;
defparam Ur0_n_2_pp.CB = 329;
defparam Ur0_n_2_pp.CC = 0;
defparam Ur0_n_2_pp.CD = 497;
defparam Ur0_n_2_pp.CE = 25;
defparam Ur0_n_2_pp.CF = 10;
wire [8:0] lut_val_0_n_3_pp;
rom_lut Ur0_n_3_pp (.addr_in( {tdl_4_n[3],tdl_2_n[3],tdl_1_n[3],tdl_0_n[3] } ), .data_out( lut_val_0_n_3_pp[8:0]) ) ;
 defparam Ur0_n_3_pp.DATA_WIDTH = 9;
defparam Ur0_n_3_pp.C0 = 0;
defparam Ur0_n_3_pp.C1 = 497;
defparam Ur0_n_3_pp.C2 = 25;
defparam Ur0_n_3_pp.C3 = 10;
defparam Ur0_n_3_pp.C4 = 193;
defparam Ur0_n_3_pp.C5 = 178;
defparam Ur0_n_3_pp.C6 = 218;
defparam Ur0_n_3_pp.C7 = 203;
defparam Ur0_n_3_pp.C8 = 319;
defparam Ur0_n_3_pp.C9 = 304;
defparam Ur0_n_3_pp.CA = 344;
defparam Ur0_n_3_pp.CB = 329;
defparam Ur0_n_3_pp.CC = 0;
defparam Ur0_n_3_pp.CD = 497;
defparam Ur0_n_3_pp.CE = 25;
defparam Ur0_n_3_pp.CF = 10;
wire [8:0] lut_val_0_n_4_pp;
rom_lut Ur0_n_4_pp (.addr_in( {tdl_4_n[4],tdl_2_n[4],tdl_1_n[4],tdl_0_n[4] } ), .data_out( lut_val_0_n_4_pp[8:0]) ) ;
 defparam Ur0_n_4_pp.DATA_WIDTH = 9;
defparam Ur0_n_4_pp.C0 = 0;
defparam Ur0_n_4_pp.C1 = 497;
defparam Ur0_n_4_pp.C2 = 25;
defparam Ur0_n_4_pp.C3 = 10;
defparam Ur0_n_4_pp.C4 = 193;
defparam Ur0_n_4_pp.C5 = 178;
defparam Ur0_n_4_pp.C6 = 218;
defparam Ur0_n_4_pp.C7 = 203;
defparam Ur0_n_4_pp.C8 = 319;
defparam Ur0_n_4_pp.C9 = 304;
defparam Ur0_n_4_pp.CA = 344;
defparam Ur0_n_4_pp.CB = 329;
defparam Ur0_n_4_pp.CC = 0;
defparam Ur0_n_4_pp.CD = 497;
defparam Ur0_n_4_pp.CE = 25;
defparam Ur0_n_4_pp.CF = 10;
wire [8:0] lut_val_0_n_5_pp;
rom_lut Ur0_n_5_pp (.addr_in( {tdl_4_n[5],tdl_2_n[5],tdl_1_n[5],tdl_0_n[5] } ), .data_out( lut_val_0_n_5_pp[8:0]) ) ;
 defparam Ur0_n_5_pp.DATA_WIDTH = 9;
defparam Ur0_n_5_pp.C0 = 0;
defparam Ur0_n_5_pp.C1 = 497;
defparam Ur0_n_5_pp.C2 = 25;
defparam Ur0_n_5_pp.C3 = 10;
defparam Ur0_n_5_pp.C4 = 193;
defparam Ur0_n_5_pp.C5 = 178;
defparam Ur0_n_5_pp.C6 = 218;
defparam Ur0_n_5_pp.C7 = 203;
defparam Ur0_n_5_pp.C8 = 319;
defparam Ur0_n_5_pp.C9 = 304;
defparam Ur0_n_5_pp.CA = 344;
defparam Ur0_n_5_pp.CB = 329;
defparam Ur0_n_5_pp.CC = 0;
defparam Ur0_n_5_pp.CD = 497;
defparam Ur0_n_5_pp.CE = 25;
defparam Ur0_n_5_pp.CF = 10;
wire [8:0] lut_val_0_n_6_pp;
rom_lut Ur0_n_6_pp (.addr_in( {tdl_4_n[6],tdl_2_n[6],tdl_1_n[6],tdl_0_n[6] } ), .data_out( lut_val_0_n_6_pp[8:0]) ) ;
 defparam Ur0_n_6_pp.DATA_WIDTH = 9;
defparam Ur0_n_6_pp.C0 = 0;
defparam Ur0_n_6_pp.C1 = 497;
defparam Ur0_n_6_pp.C2 = 25;
defparam Ur0_n_6_pp.C3 = 10;
defparam Ur0_n_6_pp.C4 = 193;
defparam Ur0_n_6_pp.C5 = 178;
defparam Ur0_n_6_pp.C6 = 218;
defparam Ur0_n_6_pp.C7 = 203;
defparam Ur0_n_6_pp.C8 = 319;
defparam Ur0_n_6_pp.C9 = 304;
defparam Ur0_n_6_pp.CA = 344;
defparam Ur0_n_6_pp.CB = 329;
defparam Ur0_n_6_pp.CC = 0;
defparam Ur0_n_6_pp.CD = 497;
defparam Ur0_n_6_pp.CE = 25;
defparam Ur0_n_6_pp.CF = 10;
wire [8:0] lut_val_0_n_7_pp;
rom_lut Ur0_n_7_pp (.addr_in( {tdl_4_n[7],tdl_2_n[7],tdl_1_n[7],tdl_0_n[7] } ), .data_out( lut_val_0_n_7_pp[8:0]) ) ;
 defparam Ur0_n_7_pp.DATA_WIDTH = 9;
defparam Ur0_n_7_pp.C0 = 0;
defparam Ur0_n_7_pp.C1 = 497;
defparam Ur0_n_7_pp.C2 = 25;
defparam Ur0_n_7_pp.C3 = 10;
defparam Ur0_n_7_pp.C4 = 193;
defparam Ur0_n_7_pp.C5 = 178;
defparam Ur0_n_7_pp.C6 = 218;
defparam Ur0_n_7_pp.C7 = 203;
defparam Ur0_n_7_pp.C8 = 319;
defparam Ur0_n_7_pp.C9 = 304;
defparam Ur0_n_7_pp.CA = 344;
defparam Ur0_n_7_pp.CB = 329;
defparam Ur0_n_7_pp.CC = 0;
defparam Ur0_n_7_pp.CD = 497;
defparam Ur0_n_7_pp.CE = 25;
defparam Ur0_n_7_pp.CF = 10;
wire [8:0] lut_val_0_n_8_pp;
rom_lut Ur0_n_8_pp (.addr_in( {tdl_4_n[8],tdl_2_n[8],tdl_1_n[8],tdl_0_n[8] } ), .data_out( lut_val_0_n_8_pp[8:0]) ) ;
 defparam Ur0_n_8_pp.DATA_WIDTH = 9;
defparam Ur0_n_8_pp.C0 = 0;
defparam Ur0_n_8_pp.C1 = 497;
defparam Ur0_n_8_pp.C2 = 25;
defparam Ur0_n_8_pp.C3 = 10;
defparam Ur0_n_8_pp.C4 = 193;
defparam Ur0_n_8_pp.C5 = 178;
defparam Ur0_n_8_pp.C6 = 218;
defparam Ur0_n_8_pp.C7 = 203;
defparam Ur0_n_8_pp.C8 = 319;
defparam Ur0_n_8_pp.C9 = 304;
defparam Ur0_n_8_pp.CA = 344;
defparam Ur0_n_8_pp.CB = 329;
defparam Ur0_n_8_pp.CC = 0;
defparam Ur0_n_8_pp.CD = 497;
defparam Ur0_n_8_pp.CE = 25;
defparam Ur0_n_8_pp.CF = 10;
wire [8:0] lut_val_0_n_9_pp;
rom_lut Ur0_n_9_pp (.addr_in( {tdl_4_n[9],tdl_2_n[9],tdl_1_n[9],tdl_0_n[9] } ), .data_out( lut_val_0_n_9_pp[8:0]) ) ;
 defparam Ur0_n_9_pp.DATA_WIDTH = 9;
defparam Ur0_n_9_pp.C0 = 0;
defparam Ur0_n_9_pp.C1 = 497;
defparam Ur0_n_9_pp.C2 = 25;
defparam Ur0_n_9_pp.C3 = 10;
defparam Ur0_n_9_pp.C4 = 193;
defparam Ur0_n_9_pp.C5 = 178;
defparam Ur0_n_9_pp.C6 = 218;
defparam Ur0_n_9_pp.C7 = 203;
defparam Ur0_n_9_pp.C8 = 319;
defparam Ur0_n_9_pp.C9 = 304;
defparam Ur0_n_9_pp.CA = 344;
defparam Ur0_n_9_pp.CB = 329;
defparam Ur0_n_9_pp.CC = 0;
defparam Ur0_n_9_pp.CD = 497;
defparam Ur0_n_9_pp.CE = 25;
defparam Ur0_n_9_pp.CF = 10;
wire [8:0] lut_val_0_n_10_pp;
rom_lut Ur0_n_10_pp (.addr_in( {tdl_4_n[10],tdl_2_n[10],tdl_1_n[10],tdl_0_n[10] } ), .data_out( lut_val_0_n_10_pp[8:0]) ) ;
 defparam Ur0_n_10_pp.DATA_WIDTH = 9;
defparam Ur0_n_10_pp.C0 = 0;
defparam Ur0_n_10_pp.C1 = 497;
defparam Ur0_n_10_pp.C2 = 25;
defparam Ur0_n_10_pp.C3 = 10;
defparam Ur0_n_10_pp.C4 = 193;
defparam Ur0_n_10_pp.C5 = 178;
defparam Ur0_n_10_pp.C6 = 218;
defparam Ur0_n_10_pp.C7 = 203;
defparam Ur0_n_10_pp.C8 = 319;
defparam Ur0_n_10_pp.C9 = 304;
defparam Ur0_n_10_pp.CA = 344;
defparam Ur0_n_10_pp.CB = 329;
defparam Ur0_n_10_pp.CC = 0;
defparam Ur0_n_10_pp.CD = 497;
defparam Ur0_n_10_pp.CE = 25;
defparam Ur0_n_10_pp.CF = 10;
wire [8:0] lut_val_0_n_11_pp;
rom_lut Ur0_n_11_pp (.addr_in( {tdl_4_n[11],tdl_2_n[11],tdl_1_n[11],tdl_0_n[11] } ), .data_out( lut_val_0_n_11_pp[8:0]) ) ;
 defparam Ur0_n_11_pp.DATA_WIDTH = 9;
defparam Ur0_n_11_pp.C0 = 0;
defparam Ur0_n_11_pp.C1 = 497;
defparam Ur0_n_11_pp.C2 = 25;
defparam Ur0_n_11_pp.C3 = 10;
defparam Ur0_n_11_pp.C4 = 193;
defparam Ur0_n_11_pp.C5 = 178;
defparam Ur0_n_11_pp.C6 = 218;
defparam Ur0_n_11_pp.C7 = 203;
defparam Ur0_n_11_pp.C8 = 319;
defparam Ur0_n_11_pp.C9 = 304;
defparam Ur0_n_11_pp.CA = 344;
defparam Ur0_n_11_pp.CB = 329;
defparam Ur0_n_11_pp.CC = 0;
defparam Ur0_n_11_pp.CD = 497;
defparam Ur0_n_11_pp.CE = 25;
defparam Ur0_n_11_pp.CF = 10;
wire [8:0] lut_val_0_n_12_pp;
rom_lut Ur0_n_12_pp (.addr_in( {tdl_4_n[12],tdl_2_n[12],tdl_1_n[12],tdl_0_n[12] } ), .data_out( lut_val_0_n_12_pp[8:0]) ) ;
 defparam Ur0_n_12_pp.DATA_WIDTH = 9;
defparam Ur0_n_12_pp.C0 = 0;
defparam Ur0_n_12_pp.C1 = 497;
defparam Ur0_n_12_pp.C2 = 25;
defparam Ur0_n_12_pp.C3 = 10;
defparam Ur0_n_12_pp.C4 = 193;
defparam Ur0_n_12_pp.C5 = 178;
defparam Ur0_n_12_pp.C6 = 218;
defparam Ur0_n_12_pp.C7 = 203;
defparam Ur0_n_12_pp.C8 = 319;
defparam Ur0_n_12_pp.C9 = 304;
defparam Ur0_n_12_pp.CA = 344;
defparam Ur0_n_12_pp.CB = 329;
defparam Ur0_n_12_pp.CC = 0;
defparam Ur0_n_12_pp.CD = 497;
defparam Ur0_n_12_pp.CE = 25;
defparam Ur0_n_12_pp.CF = 10;
wire [8:0] lut_val_0_n_13_pp;
rom_lut Ur0_n_13_pp (.addr_in( {tdl_4_n[13],tdl_2_n[13],tdl_1_n[13],tdl_0_n[13] } ), .data_out( lut_val_0_n_13_pp[8:0]) ) ;
 defparam Ur0_n_13_pp.DATA_WIDTH = 9;
defparam Ur0_n_13_pp.C0 = 0;
defparam Ur0_n_13_pp.C1 = 497;
defparam Ur0_n_13_pp.C2 = 25;
defparam Ur0_n_13_pp.C3 = 10;
defparam Ur0_n_13_pp.C4 = 193;
defparam Ur0_n_13_pp.C5 = 178;
defparam Ur0_n_13_pp.C6 = 218;
defparam Ur0_n_13_pp.C7 = 203;
defparam Ur0_n_13_pp.C8 = 319;
defparam Ur0_n_13_pp.C9 = 304;
defparam Ur0_n_13_pp.CA = 344;
defparam Ur0_n_13_pp.CB = 329;
defparam Ur0_n_13_pp.CC = 0;
defparam Ur0_n_13_pp.CD = 497;
defparam Ur0_n_13_pp.CE = 25;
defparam Ur0_n_13_pp.CF = 10;
wire [8:0] lut_val_0_n_14_pp;
rom_lut Ur0_n_14_pp (.addr_in( {tdl_4_n[14],tdl_2_n[14],tdl_1_n[14],tdl_0_n[14] } ), .data_out( lut_val_0_n_14_pp[8:0]) ) ;
 defparam Ur0_n_14_pp.DATA_WIDTH = 9;
defparam Ur0_n_14_pp.C0 = 0;
defparam Ur0_n_14_pp.C1 = 497;
defparam Ur0_n_14_pp.C2 = 25;
defparam Ur0_n_14_pp.C3 = 10;
defparam Ur0_n_14_pp.C4 = 193;
defparam Ur0_n_14_pp.C5 = 178;
defparam Ur0_n_14_pp.C6 = 218;
defparam Ur0_n_14_pp.C7 = 203;
defparam Ur0_n_14_pp.C8 = 319;
defparam Ur0_n_14_pp.C9 = 304;
defparam Ur0_n_14_pp.CA = 344;
defparam Ur0_n_14_pp.CB = 329;
defparam Ur0_n_14_pp.CC = 0;
defparam Ur0_n_14_pp.CD = 497;
defparam Ur0_n_14_pp.CE = 25;
defparam Ur0_n_14_pp.CF = 10;
wire [8:0] lut_val_0_n_15_pp;
rom_lut Ur0_n_15_pp (.addr_in( {tdl_4_n[15],tdl_2_n[15],tdl_1_n[15],tdl_0_n[15] } ), .data_out( lut_val_0_n_15_pp[8:0]) ) ;
 defparam Ur0_n_15_pp.DATA_WIDTH = 9;
defparam Ur0_n_15_pp.C0 = 0;
defparam Ur0_n_15_pp.C1 = 15;
defparam Ur0_n_15_pp.C2 = 487;
defparam Ur0_n_15_pp.C3 = 502;
defparam Ur0_n_15_pp.C4 = 319;
defparam Ur0_n_15_pp.C5 = 334;
defparam Ur0_n_15_pp.C6 = 294;
defparam Ur0_n_15_pp.C7 = 309;
defparam Ur0_n_15_pp.C8 = 193;
defparam Ur0_n_15_pp.C9 = 208;
defparam Ur0_n_15_pp.CA = 168;
defparam Ur0_n_15_pp.CB = 183;
defparam Ur0_n_15_pp.CC = 0;
defparam Ur0_n_15_pp.CD = 15;
defparam Ur0_n_15_pp.CE = 487;
defparam Ur0_n_15_pp.CF = 502;
wire [8:0] lut_val_1_n_0_pp;
rom_lut Ur1_n_0_pp (.addr_in( {addr_low,addr_low,tdl_6_n[0],tdl_5_n[0] } ), .data_out( lut_val_1_n_0_pp[5:0]) ) ;
 defparam Ur1_n_0_pp.DATA_WIDTH = 6;
defparam Ur1_n_0_pp.C0 = 0;
defparam Ur1_n_0_pp.C1 = 39;
defparam Ur1_n_0_pp.C2 = 15;
defparam Ur1_n_0_pp.C3 = 54;
defparam Ur1_n_0_pp.C4 = 0;
defparam Ur1_n_0_pp.C5 = 39;
defparam Ur1_n_0_pp.C6 = 15;
defparam Ur1_n_0_pp.C7 = 54;
defparam Ur1_n_0_pp.C8 = 0;
defparam Ur1_n_0_pp.C9 = 39;
defparam Ur1_n_0_pp.CA = 15;
defparam Ur1_n_0_pp.CB = 54;
defparam Ur1_n_0_pp.CC = 0;
defparam Ur1_n_0_pp.CD = 39;
defparam Ur1_n_0_pp.CE = 15;
defparam Ur1_n_0_pp.CF = 54;
assign lut_val_1_n_0_pp[8] = lut_val_1_n_0_pp[5];
assign lut_val_1_n_0_pp[7] = lut_val_1_n_0_pp[5];
assign lut_val_1_n_0_pp[6] = lut_val_1_n_0_pp[5];
wire [8:0] lut_val_1_n_1_pp;
rom_lut Ur1_n_1_pp (.addr_in( {addr_low,addr_low,tdl_6_n[1],tdl_5_n[1] } ), .data_out( lut_val_1_n_1_pp[5:0]) ) ;
 defparam Ur1_n_1_pp.DATA_WIDTH = 6;
defparam Ur1_n_1_pp.C0 = 0;
defparam Ur1_n_1_pp.C1 = 39;
defparam Ur1_n_1_pp.C2 = 15;
defparam Ur1_n_1_pp.C3 = 54;
defparam Ur1_n_1_pp.C4 = 0;
defparam Ur1_n_1_pp.C5 = 39;
defparam Ur1_n_1_pp.C6 = 15;
defparam Ur1_n_1_pp.C7 = 54;
defparam Ur1_n_1_pp.C8 = 0;
defparam Ur1_n_1_pp.C9 = 39;
defparam Ur1_n_1_pp.CA = 15;
defparam Ur1_n_1_pp.CB = 54;
defparam Ur1_n_1_pp.CC = 0;
defparam Ur1_n_1_pp.CD = 39;
defparam Ur1_n_1_pp.CE = 15;
defparam Ur1_n_1_pp.CF = 54;
assign lut_val_1_n_1_pp[8] = lut_val_1_n_1_pp[5];
assign lut_val_1_n_1_pp[7] = lut_val_1_n_1_pp[5];
assign lut_val_1_n_1_pp[6] = lut_val_1_n_1_pp[5];
wire [8:0] lut_val_1_n_2_pp;
rom_lut Ur1_n_2_pp (.addr_in( {addr_low,addr_low,tdl_6_n[2],tdl_5_n[2] } ), .data_out( lut_val_1_n_2_pp[5:0]) ) ;
 defparam Ur1_n_2_pp.DATA_WIDTH = 6;
defparam Ur1_n_2_pp.C0 = 0;
defparam Ur1_n_2_pp.C1 = 39;
defparam Ur1_n_2_pp.C2 = 15;
defparam Ur1_n_2_pp.C3 = 54;
defparam Ur1_n_2_pp.C4 = 0;
defparam Ur1_n_2_pp.C5 = 39;
defparam Ur1_n_2_pp.C6 = 15;
defparam Ur1_n_2_pp.C7 = 54;
defparam Ur1_n_2_pp.C8 = 0;
defparam Ur1_n_2_pp.C9 = 39;
defparam Ur1_n_2_pp.CA = 15;
defparam Ur1_n_2_pp.CB = 54;
defparam Ur1_n_2_pp.CC = 0;
defparam Ur1_n_2_pp.CD = 39;
defparam Ur1_n_2_pp.CE = 15;
defparam Ur1_n_2_pp.CF = 54;
assign lut_val_1_n_2_pp[8] = lut_val_1_n_2_pp[5];
assign lut_val_1_n_2_pp[7] = lut_val_1_n_2_pp[5];
assign lut_val_1_n_2_pp[6] = lut_val_1_n_2_pp[5];
wire [8:0] lut_val_1_n_3_pp;
rom_lut Ur1_n_3_pp (.addr_in( {addr_low,addr_low,tdl_6_n[3],tdl_5_n[3] } ), .data_out( lut_val_1_n_3_pp[5:0]) ) ;
 defparam Ur1_n_3_pp.DATA_WIDTH = 6;
defparam Ur1_n_3_pp.C0 = 0;
defparam Ur1_n_3_pp.C1 = 39;
defparam Ur1_n_3_pp.C2 = 15;
defparam Ur1_n_3_pp.C3 = 54;
defparam Ur1_n_3_pp.C4 = 0;
defparam Ur1_n_3_pp.C5 = 39;
defparam Ur1_n_3_pp.C6 = 15;
defparam Ur1_n_3_pp.C7 = 54;
defparam Ur1_n_3_pp.C8 = 0;
defparam Ur1_n_3_pp.C9 = 39;
defparam Ur1_n_3_pp.CA = 15;
defparam Ur1_n_3_pp.CB = 54;
defparam Ur1_n_3_pp.CC = 0;
defparam Ur1_n_3_pp.CD = 39;
defparam Ur1_n_3_pp.CE = 15;
defparam Ur1_n_3_pp.CF = 54;
assign lut_val_1_n_3_pp[8] = lut_val_1_n_3_pp[5];
assign lut_val_1_n_3_pp[7] = lut_val_1_n_3_pp[5];
assign lut_val_1_n_3_pp[6] = lut_val_1_n_3_pp[5];
wire [8:0] lut_val_1_n_4_pp;
rom_lut Ur1_n_4_pp (.addr_in( {addr_low,addr_low,tdl_6_n[4],tdl_5_n[4] } ), .data_out( lut_val_1_n_4_pp[5:0]) ) ;
 defparam Ur1_n_4_pp.DATA_WIDTH = 6;
defparam Ur1_n_4_pp.C0 = 0;
defparam Ur1_n_4_pp.C1 = 39;
defparam Ur1_n_4_pp.C2 = 15;
defparam Ur1_n_4_pp.C3 = 54;
defparam Ur1_n_4_pp.C4 = 0;
defparam Ur1_n_4_pp.C5 = 39;
defparam Ur1_n_4_pp.C6 = 15;
defparam Ur1_n_4_pp.C7 = 54;
defparam Ur1_n_4_pp.C8 = 0;
defparam Ur1_n_4_pp.C9 = 39;
defparam Ur1_n_4_pp.CA = 15;
defparam Ur1_n_4_pp.CB = 54;
defparam Ur1_n_4_pp.CC = 0;
defparam Ur1_n_4_pp.CD = 39;
defparam Ur1_n_4_pp.CE = 15;
defparam Ur1_n_4_pp.CF = 54;
assign lut_val_1_n_4_pp[8] = lut_val_1_n_4_pp[5];
assign lut_val_1_n_4_pp[7] = lut_val_1_n_4_pp[5];
assign lut_val_1_n_4_pp[6] = lut_val_1_n_4_pp[5];
wire [8:0] lut_val_1_n_5_pp;
rom_lut Ur1_n_5_pp (.addr_in( {addr_low,addr_low,tdl_6_n[5],tdl_5_n[5] } ), .data_out( lut_val_1_n_5_pp[5:0]) ) ;
 defparam Ur1_n_5_pp.DATA_WIDTH = 6;
defparam Ur1_n_5_pp.C0 = 0;
defparam Ur1_n_5_pp.C1 = 39;
defparam Ur1_n_5_pp.C2 = 15;
defparam Ur1_n_5_pp.C3 = 54;
defparam Ur1_n_5_pp.C4 = 0;
defparam Ur1_n_5_pp.C5 = 39;
defparam Ur1_n_5_pp.C6 = 15;
defparam Ur1_n_5_pp.C7 = 54;
defparam Ur1_n_5_pp.C8 = 0;
defparam Ur1_n_5_pp.C9 = 39;
defparam Ur1_n_5_pp.CA = 15;
defparam Ur1_n_5_pp.CB = 54;
defparam Ur1_n_5_pp.CC = 0;
defparam Ur1_n_5_pp.CD = 39;
defparam Ur1_n_5_pp.CE = 15;
defparam Ur1_n_5_pp.CF = 54;
assign lut_val_1_n_5_pp[8] = lut_val_1_n_5_pp[5];
assign lut_val_1_n_5_pp[7] = lut_val_1_n_5_pp[5];
assign lut_val_1_n_5_pp[6] = lut_val_1_n_5_pp[5];
wire [8:0] lut_val_1_n_6_pp;
rom_lut Ur1_n_6_pp (.addr_in( {addr_low,addr_low,tdl_6_n[6],tdl_5_n[6] } ), .data_out( lut_val_1_n_6_pp[5:0]) ) ;
 defparam Ur1_n_6_pp.DATA_WIDTH = 6;
defparam Ur1_n_6_pp.C0 = 0;
defparam Ur1_n_6_pp.C1 = 39;
defparam Ur1_n_6_pp.C2 = 15;
defparam Ur1_n_6_pp.C3 = 54;
defparam Ur1_n_6_pp.C4 = 0;
defparam Ur1_n_6_pp.C5 = 39;
defparam Ur1_n_6_pp.C6 = 15;
defparam Ur1_n_6_pp.C7 = 54;
defparam Ur1_n_6_pp.C8 = 0;
defparam Ur1_n_6_pp.C9 = 39;
defparam Ur1_n_6_pp.CA = 15;
defparam Ur1_n_6_pp.CB = 54;
defparam Ur1_n_6_pp.CC = 0;
defparam Ur1_n_6_pp.CD = 39;
defparam Ur1_n_6_pp.CE = 15;
defparam Ur1_n_6_pp.CF = 54;
assign lut_val_1_n_6_pp[8] = lut_val_1_n_6_pp[5];
assign lut_val_1_n_6_pp[7] = lut_val_1_n_6_pp[5];
assign lut_val_1_n_6_pp[6] = lut_val_1_n_6_pp[5];
wire [8:0] lut_val_1_n_7_pp;
rom_lut Ur1_n_7_pp (.addr_in( {addr_low,addr_low,tdl_6_n[7],tdl_5_n[7] } ), .data_out( lut_val_1_n_7_pp[5:0]) ) ;
 defparam Ur1_n_7_pp.DATA_WIDTH = 6;
defparam Ur1_n_7_pp.C0 = 0;
defparam Ur1_n_7_pp.C1 = 39;
defparam Ur1_n_7_pp.C2 = 15;
defparam Ur1_n_7_pp.C3 = 54;
defparam Ur1_n_7_pp.C4 = 0;
defparam Ur1_n_7_pp.C5 = 39;
defparam Ur1_n_7_pp.C6 = 15;
defparam Ur1_n_7_pp.C7 = 54;
defparam Ur1_n_7_pp.C8 = 0;
defparam Ur1_n_7_pp.C9 = 39;
defparam Ur1_n_7_pp.CA = 15;
defparam Ur1_n_7_pp.CB = 54;
defparam Ur1_n_7_pp.CC = 0;
defparam Ur1_n_7_pp.CD = 39;
defparam Ur1_n_7_pp.CE = 15;
defparam Ur1_n_7_pp.CF = 54;
assign lut_val_1_n_7_pp[8] = lut_val_1_n_7_pp[5];
assign lut_val_1_n_7_pp[7] = lut_val_1_n_7_pp[5];
assign lut_val_1_n_7_pp[6] = lut_val_1_n_7_pp[5];
wire [8:0] lut_val_1_n_8_pp;
rom_lut Ur1_n_8_pp (.addr_in( {addr_low,addr_low,tdl_6_n[8],tdl_5_n[8] } ), .data_out( lut_val_1_n_8_pp[5:0]) ) ;
 defparam Ur1_n_8_pp.DATA_WIDTH = 6;
defparam Ur1_n_8_pp.C0 = 0;
defparam Ur1_n_8_pp.C1 = 39;
defparam Ur1_n_8_pp.C2 = 15;
defparam Ur1_n_8_pp.C3 = 54;
defparam Ur1_n_8_pp.C4 = 0;
defparam Ur1_n_8_pp.C5 = 39;
defparam Ur1_n_8_pp.C6 = 15;
defparam Ur1_n_8_pp.C7 = 54;
defparam Ur1_n_8_pp.C8 = 0;
defparam Ur1_n_8_pp.C9 = 39;
defparam Ur1_n_8_pp.CA = 15;
defparam Ur1_n_8_pp.CB = 54;
defparam Ur1_n_8_pp.CC = 0;
defparam Ur1_n_8_pp.CD = 39;
defparam Ur1_n_8_pp.CE = 15;
defparam Ur1_n_8_pp.CF = 54;
assign lut_val_1_n_8_pp[8] = lut_val_1_n_8_pp[5];
assign lut_val_1_n_8_pp[7] = lut_val_1_n_8_pp[5];
assign lut_val_1_n_8_pp[6] = lut_val_1_n_8_pp[5];
wire [8:0] lut_val_1_n_9_pp;
rom_lut Ur1_n_9_pp (.addr_in( {addr_low,addr_low,tdl_6_n[9],tdl_5_n[9] } ), .data_out( lut_val_1_n_9_pp[5:0]) ) ;
 defparam Ur1_n_9_pp.DATA_WIDTH = 6;
defparam Ur1_n_9_pp.C0 = 0;
defparam Ur1_n_9_pp.C1 = 39;
defparam Ur1_n_9_pp.C2 = 15;
defparam Ur1_n_9_pp.C3 = 54;
defparam Ur1_n_9_pp.C4 = 0;
defparam Ur1_n_9_pp.C5 = 39;
defparam Ur1_n_9_pp.C6 = 15;
defparam Ur1_n_9_pp.C7 = 54;
defparam Ur1_n_9_pp.C8 = 0;
defparam Ur1_n_9_pp.C9 = 39;
defparam Ur1_n_9_pp.CA = 15;
defparam Ur1_n_9_pp.CB = 54;
defparam Ur1_n_9_pp.CC = 0;
defparam Ur1_n_9_pp.CD = 39;
defparam Ur1_n_9_pp.CE = 15;
defparam Ur1_n_9_pp.CF = 54;
assign lut_val_1_n_9_pp[8] = lut_val_1_n_9_pp[5];
assign lut_val_1_n_9_pp[7] = lut_val_1_n_9_pp[5];
assign lut_val_1_n_9_pp[6] = lut_val_1_n_9_pp[5];
wire [8:0] lut_val_1_n_10_pp;
rom_lut Ur1_n_10_pp (.addr_in( {addr_low,addr_low,tdl_6_n[10],tdl_5_n[10] } ), .data_out( lut_val_1_n_10_pp[5:0]) ) ;
 defparam Ur1_n_10_pp.DATA_WIDTH = 6;
defparam Ur1_n_10_pp.C0 = 0;
defparam Ur1_n_10_pp.C1 = 39;
defparam Ur1_n_10_pp.C2 = 15;
defparam Ur1_n_10_pp.C3 = 54;
defparam Ur1_n_10_pp.C4 = 0;
defparam Ur1_n_10_pp.C5 = 39;
defparam Ur1_n_10_pp.C6 = 15;
defparam Ur1_n_10_pp.C7 = 54;
defparam Ur1_n_10_pp.C8 = 0;
defparam Ur1_n_10_pp.C9 = 39;
defparam Ur1_n_10_pp.CA = 15;
defparam Ur1_n_10_pp.CB = 54;
defparam Ur1_n_10_pp.CC = 0;
defparam Ur1_n_10_pp.CD = 39;
defparam Ur1_n_10_pp.CE = 15;
defparam Ur1_n_10_pp.CF = 54;
assign lut_val_1_n_10_pp[8] = lut_val_1_n_10_pp[5];
assign lut_val_1_n_10_pp[7] = lut_val_1_n_10_pp[5];
assign lut_val_1_n_10_pp[6] = lut_val_1_n_10_pp[5];
wire [8:0] lut_val_1_n_11_pp;
rom_lut Ur1_n_11_pp (.addr_in( {addr_low,addr_low,tdl_6_n[11],tdl_5_n[11] } ), .data_out( lut_val_1_n_11_pp[5:0]) ) ;
 defparam Ur1_n_11_pp.DATA_WIDTH = 6;
defparam Ur1_n_11_pp.C0 = 0;
defparam Ur1_n_11_pp.C1 = 39;
defparam Ur1_n_11_pp.C2 = 15;
defparam Ur1_n_11_pp.C3 = 54;
defparam Ur1_n_11_pp.C4 = 0;
defparam Ur1_n_11_pp.C5 = 39;
defparam Ur1_n_11_pp.C6 = 15;
defparam Ur1_n_11_pp.C7 = 54;
defparam Ur1_n_11_pp.C8 = 0;
defparam Ur1_n_11_pp.C9 = 39;
defparam Ur1_n_11_pp.CA = 15;
defparam Ur1_n_11_pp.CB = 54;
defparam Ur1_n_11_pp.CC = 0;
defparam Ur1_n_11_pp.CD = 39;
defparam Ur1_n_11_pp.CE = 15;
defparam Ur1_n_11_pp.CF = 54;
assign lut_val_1_n_11_pp[8] = lut_val_1_n_11_pp[5];
assign lut_val_1_n_11_pp[7] = lut_val_1_n_11_pp[5];
assign lut_val_1_n_11_pp[6] = lut_val_1_n_11_pp[5];
wire [8:0] lut_val_1_n_12_pp;
rom_lut Ur1_n_12_pp (.addr_in( {addr_low,addr_low,tdl_6_n[12],tdl_5_n[12] } ), .data_out( lut_val_1_n_12_pp[5:0]) ) ;
 defparam Ur1_n_12_pp.DATA_WIDTH = 6;
defparam Ur1_n_12_pp.C0 = 0;
defparam Ur1_n_12_pp.C1 = 39;
defparam Ur1_n_12_pp.C2 = 15;
defparam Ur1_n_12_pp.C3 = 54;
defparam Ur1_n_12_pp.C4 = 0;
defparam Ur1_n_12_pp.C5 = 39;
defparam Ur1_n_12_pp.C6 = 15;
defparam Ur1_n_12_pp.C7 = 54;
defparam Ur1_n_12_pp.C8 = 0;
defparam Ur1_n_12_pp.C9 = 39;
defparam Ur1_n_12_pp.CA = 15;
defparam Ur1_n_12_pp.CB = 54;
defparam Ur1_n_12_pp.CC = 0;
defparam Ur1_n_12_pp.CD = 39;
defparam Ur1_n_12_pp.CE = 15;
defparam Ur1_n_12_pp.CF = 54;
assign lut_val_1_n_12_pp[8] = lut_val_1_n_12_pp[5];
assign lut_val_1_n_12_pp[7] = lut_val_1_n_12_pp[5];
assign lut_val_1_n_12_pp[6] = lut_val_1_n_12_pp[5];
wire [8:0] lut_val_1_n_13_pp;
rom_lut Ur1_n_13_pp (.addr_in( {addr_low,addr_low,tdl_6_n[13],tdl_5_n[13] } ), .data_out( lut_val_1_n_13_pp[5:0]) ) ;
 defparam Ur1_n_13_pp.DATA_WIDTH = 6;
defparam Ur1_n_13_pp.C0 = 0;
defparam Ur1_n_13_pp.C1 = 39;
defparam Ur1_n_13_pp.C2 = 15;
defparam Ur1_n_13_pp.C3 = 54;
defparam Ur1_n_13_pp.C4 = 0;
defparam Ur1_n_13_pp.C5 = 39;
defparam Ur1_n_13_pp.C6 = 15;
defparam Ur1_n_13_pp.C7 = 54;
defparam Ur1_n_13_pp.C8 = 0;
defparam Ur1_n_13_pp.C9 = 39;
defparam Ur1_n_13_pp.CA = 15;
defparam Ur1_n_13_pp.CB = 54;
defparam Ur1_n_13_pp.CC = 0;
defparam Ur1_n_13_pp.CD = 39;
defparam Ur1_n_13_pp.CE = 15;
defparam Ur1_n_13_pp.CF = 54;
assign lut_val_1_n_13_pp[8] = lut_val_1_n_13_pp[5];
assign lut_val_1_n_13_pp[7] = lut_val_1_n_13_pp[5];
assign lut_val_1_n_13_pp[6] = lut_val_1_n_13_pp[5];
wire [8:0] lut_val_1_n_14_pp;
rom_lut Ur1_n_14_pp (.addr_in( {addr_low,addr_low,tdl_6_n[14],tdl_5_n[14] } ), .data_out( lut_val_1_n_14_pp[5:0]) ) ;
 defparam Ur1_n_14_pp.DATA_WIDTH = 6;
defparam Ur1_n_14_pp.C0 = 0;
defparam Ur1_n_14_pp.C1 = 39;
defparam Ur1_n_14_pp.C2 = 15;
defparam Ur1_n_14_pp.C3 = 54;
defparam Ur1_n_14_pp.C4 = 0;
defparam Ur1_n_14_pp.C5 = 39;
defparam Ur1_n_14_pp.C6 = 15;
defparam Ur1_n_14_pp.C7 = 54;
defparam Ur1_n_14_pp.C8 = 0;
defparam Ur1_n_14_pp.C9 = 39;
defparam Ur1_n_14_pp.CA = 15;
defparam Ur1_n_14_pp.CB = 54;
defparam Ur1_n_14_pp.CC = 0;
defparam Ur1_n_14_pp.CD = 39;
defparam Ur1_n_14_pp.CE = 15;
defparam Ur1_n_14_pp.CF = 54;
assign lut_val_1_n_14_pp[8] = lut_val_1_n_14_pp[5];
assign lut_val_1_n_14_pp[7] = lut_val_1_n_14_pp[5];
assign lut_val_1_n_14_pp[6] = lut_val_1_n_14_pp[5];
wire [8:0] lut_val_1_n_15_pp;
rom_lut Ur1_n_15_pp (.addr_in( {addr_low,addr_low,tdl_6_n[15],tdl_5_n[15] } ), .data_out( lut_val_1_n_15_pp[5:0]) ) ;
 defparam Ur1_n_15_pp.DATA_WIDTH = 6;
defparam Ur1_n_15_pp.C0 = 0;
defparam Ur1_n_15_pp.C1 = 25;
defparam Ur1_n_15_pp.C2 = 49;
defparam Ur1_n_15_pp.C3 = 10;
defparam Ur1_n_15_pp.C4 = 0;
defparam Ur1_n_15_pp.C5 = 25;
defparam Ur1_n_15_pp.C6 = 49;
defparam Ur1_n_15_pp.C7 = 10;
defparam Ur1_n_15_pp.C8 = 0;
defparam Ur1_n_15_pp.C9 = 25;
defparam Ur1_n_15_pp.CA = 49;
defparam Ur1_n_15_pp.CB = 10;
defparam Ur1_n_15_pp.CC = 0;
defparam Ur1_n_15_pp.CD = 25;
defparam Ur1_n_15_pp.CE = 49;
defparam Ur1_n_15_pp.CF = 10;
assign lut_val_1_n_15_pp[8] = lut_val_1_n_15_pp[5];
assign lut_val_1_n_15_pp[7] = lut_val_1_n_15_pp[5];
assign lut_val_1_n_15_pp[6] = lut_val_1_n_15_pp[5];


// ---- partial product adder tree ----

wire [23:0] lut_0_bit_0_fill;
wire [23:0] lut_0_bit_1_fill;
wire [23:0] lut_0_bit_2_fill;
wire [23:0] lut_0_bit_3_fill;
wire [23:0] lut_0_bit_4_fill;
wire [23:0] lut_0_bit_5_fill;
wire [23:0] lut_0_bit_6_fill;
wire [23:0] lut_0_bit_7_fill;
wire [23:0] lut_0_bit_8_fill;
wire [23:0] lut_0_bit_9_fill;
wire [23:0] lut_0_bit_10_fill;
wire [23:0] lut_0_bit_11_fill;
wire [23:0] lut_0_bit_12_fill;
wire [23:0] lut_0_bit_13_fill;
wire [23:0] lut_0_bit_14_fill;
wire [23:0] lut_0_bit_15_fill;
assign lut_0_bit_0_fill = {lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8], lut_val_0_n_0_pp[8],  lut_val_0_n_0_pp };
assign lut_0_bit_1_fill = {lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8], lut_val_0_n_1_pp[8],  lut_val_0_n_1_pp, 1'd0 };
assign lut_0_bit_2_fill = {lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8], lut_val_0_n_2_pp[8],  lut_val_0_n_2_pp, 2'd0 };
assign lut_0_bit_3_fill = {lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8], lut_val_0_n_3_pp[8],  lut_val_0_n_3_pp, 3'd0 };
assign lut_0_bit_4_fill = {lut_val_0_n_4_pp[8], lut_val_0_n_4_pp[8], lut_val_0_n_4_pp[8], lut_val_0_n_4_pp[8], lut_val_0_n_4_pp[8], lut_val_0_n_4_pp[8], lut_val_0_n_4_pp[8], lut_val_0_n_4_pp[8], lut_val_0_n_4_pp[8], lut_val_0_n_4_pp[8], lut_val_0_n_4_pp[8],  lut_val_0_n_4_pp, 4'd0 };
assign lut_0_bit_5_fill = {lut_val_0_n_5_pp[8], lut_val_0_n_5_pp[8], lut_val_0_n_5_pp[8], lut_val_0_n_5_pp[8], lut_val_0_n_5_pp[8], lut_val_0_n_5_pp[8], lut_val_0_n_5_pp[8], lut_val_0_n_5_pp[8], lut_val_0_n_5_pp[8], lut_val_0_n_5_pp[8],  lut_val_0_n_5_pp, 5'd0 };
assign lut_0_bit_6_fill = {lut_val_0_n_6_pp[8], lut_val_0_n_6_pp[8], lut_val_0_n_6_pp[8], lut_val_0_n_6_pp[8], lut_val_0_n_6_pp[8], lut_val_0_n_6_pp[8], lut_val_0_n_6_pp[8], lut_val_0_n_6_pp[8], lut_val_0_n_6_pp[8],  lut_val_0_n_6_pp, 6'd0 };
assign lut_0_bit_7_fill = {lut_val_0_n_7_pp[8], lut_val_0_n_7_pp[8], lut_val_0_n_7_pp[8], lut_val_0_n_7_pp[8], lut_val_0_n_7_pp[8], lut_val_0_n_7_pp[8], lut_val_0_n_7_pp[8], lut_val_0_n_7_pp[8],  lut_val_0_n_7_pp, 7'd0 };
assign lut_0_bit_8_fill = {lut_val_0_n_8_pp[8], lut_val_0_n_8_pp[8], lut_val_0_n_8_pp[8], lut_val_0_n_8_pp[8], lut_val_0_n_8_pp[8], lut_val_0_n_8_pp[8], lut_val_0_n_8_pp[8],  lut_val_0_n_8_pp, 8'd0 };
assign lut_0_bit_9_fill = {lut_val_0_n_9_pp[8], lut_val_0_n_9_pp[8], lut_val_0_n_9_pp[8], lut_val_0_n_9_pp[8], lut_val_0_n_9_pp[8], lut_val_0_n_9_pp[8],  lut_val_0_n_9_pp, 9'd0 };
assign lut_0_bit_10_fill = {lut_val_0_n_10_pp[8], lut_val_0_n_10_pp[8], lut_val_0_n_10_pp[8], lut_val_0_n_10_pp[8], lut_val_0_n_10_pp[8],  lut_val_0_n_10_pp, 10'd0 };
assign lut_0_bit_11_fill = {lut_val_0_n_11_pp[8], lut_val_0_n_11_pp[8], lut_val_0_n_11_pp[8], lut_val_0_n_11_pp[8],  lut_val_0_n_11_pp, 11'd0 };
assign lut_0_bit_12_fill = {lut_val_0_n_12_pp[8], lut_val_0_n_12_pp[8], lut_val_0_n_12_pp[8],  lut_val_0_n_12_pp, 12'd0 };
assign lut_0_bit_13_fill = {lut_val_0_n_13_pp[8], lut_val_0_n_13_pp[8],  lut_val_0_n_13_pp, 13'd0 };
assign lut_0_bit_14_fill = {lut_val_0_n_14_pp[8],  lut_val_0_n_14_pp, 14'd0 };
assign lut_0_bit_15_fill = { lut_val_0_n_15_pp, 15'd0 };
wire [24:0] tree_0_pp_l_0_n_0_n;
sadd_lpm Uadd_0_lut_l_0_n_0_n (.clk(clk), .ain(lut_0_bit_0_fill), .bin(lut_0_bit_1_fill), .res(tree_0_pp_l_0_n_0_n) );
defparam Uadd_0_lut_l_0_n_0_n.IN_WIDTH = 24;
defparam Uadd_0_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [24:0] tree_0_pp_l_0_n_1_n;
sadd_lpm Uadd_0_lut_l_0_n_1_n (.clk(clk), .ain(lut_0_bit_2_fill), .bin(lut_0_bit_3_fill), .res(tree_0_pp_l_0_n_1_n) );
defparam Uadd_0_lut_l_0_n_1_n.IN_WIDTH = 24;
defparam Uadd_0_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [24:0] tree_0_pp_l_0_n_2_n;
sadd_lpm Uadd_0_lut_l_0_n_2_n (.clk(clk), .ain(lut_0_bit_4_fill), .bin(lut_0_bit_5_fill), .res(tree_0_pp_l_0_n_2_n) );
defparam Uadd_0_lut_l_0_n_2_n.IN_WIDTH = 24;
defparam Uadd_0_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [24:0] tree_0_pp_l_0_n_3_n;
sadd_lpm Uadd_0_lut_l_0_n_3_n (.clk(clk), .ain(lut_0_bit_6_fill), .bin(lut_0_bit_7_fill), .res(tree_0_pp_l_0_n_3_n) );
defparam Uadd_0_lut_l_0_n_3_n.IN_WIDTH = 24;
defparam Uadd_0_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [24:0] tree_0_pp_l_0_n_4_n;
sadd_lpm Uadd_0_lut_l_0_n_4_n (.clk(clk), .ain(lut_0_bit_8_fill), .bin(lut_0_bit_9_fill), .res(tree_0_pp_l_0_n_4_n) );
defparam Uadd_0_lut_l_0_n_4_n.IN_WIDTH = 24;
defparam Uadd_0_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [24:0] tree_0_pp_l_0_n_5_n;
sadd_lpm Uadd_0_lut_l_0_n_5_n (.clk(clk), .ain(lut_0_bit_10_fill), .bin(lut_0_bit_11_fill), .res(tree_0_pp_l_0_n_5_n) );
defparam Uadd_0_lut_l_0_n_5_n.IN_WIDTH = 24;
defparam Uadd_0_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [24:0] tree_0_pp_l_0_n_6_n;
sadd_lpm Uadd_0_lut_l_0_n_6_n (.clk(clk), .ain(lut_0_bit_12_fill), .bin(lut_0_bit_13_fill), .res(tree_0_pp_l_0_n_6_n) );
defparam Uadd_0_lut_l_0_n_6_n.IN_WIDTH = 24;
defparam Uadd_0_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [24:0] tree_0_pp_l_0_n_7_n;
sadd_lpm Uadd_0_lut_l_0_n_7_n (.clk(clk), .ain(lut_0_bit_14_fill), .bin(lut_0_bit_15_fill), .res(tree_0_pp_l_0_n_7_n) );
defparam Uadd_0_lut_l_0_n_7_n.IN_WIDTH = 24;
defparam Uadd_0_lut_l_0_n_7_n.PIPE_DEPTH = 1;

wire [25:0] tree_0_pp_l_1_n_0_n;
sadd_lpm Uadd_0_lut_l_1_n_0_n (.clk(clk), .ain(tree_0_pp_l_0_n_0_n), .bin(tree_0_pp_l_0_n_1_n), .res(tree_0_pp_l_1_n_0_n) );
defparam Uadd_0_lut_l_1_n_0_n.IN_WIDTH = 25;
defparam Uadd_0_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [25:0] tree_0_pp_l_1_n_1_n;
sadd_lpm Uadd_0_lut_l_1_n_1_n (.clk(clk), .ain(tree_0_pp_l_0_n_2_n), .bin(tree_0_pp_l_0_n_3_n), .res(tree_0_pp_l_1_n_1_n) );
defparam Uadd_0_lut_l_1_n_1_n.IN_WIDTH = 25;
defparam Uadd_0_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [25:0] tree_0_pp_l_1_n_2_n;
sadd_lpm Uadd_0_lut_l_1_n_2_n (.clk(clk), .ain(tree_0_pp_l_0_n_4_n), .bin(tree_0_pp_l_0_n_5_n), .res(tree_0_pp_l_1_n_2_n) );
defparam Uadd_0_lut_l_1_n_2_n.IN_WIDTH = 25;
defparam Uadd_0_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [25:0] tree_0_pp_l_1_n_3_n;
sadd_lpm Uadd_0_lut_l_1_n_3_n (.clk(clk), .ain(tree_0_pp_l_0_n_6_n), .bin(tree_0_pp_l_0_n_7_n), .res(tree_0_pp_l_1_n_3_n) );
defparam Uadd_0_lut_l_1_n_3_n.IN_WIDTH = 25;
defparam Uadd_0_lut_l_1_n_3_n.PIPE_DEPTH = 1;

wire [26:0] tree_0_pp_l_2_n_0_n;
sadd_lpm Uadd_0_lut_l_2_n_0_n (.clk(clk), .ain(tree_0_pp_l_1_n_0_n), .bin(tree_0_pp_l_1_n_1_n), .res(tree_0_pp_l_2_n_0_n) );
defparam Uadd_0_lut_l_2_n_0_n.IN_WIDTH = 26;
defparam Uadd_0_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [26:0] tree_0_pp_l_2_n_1_n;
sadd_lpm Uadd_0_lut_l_2_n_1_n (.clk(clk), .ain(tree_0_pp_l_1_n_2_n), .bin(tree_0_pp_l_1_n_3_n), .res(tree_0_pp_l_2_n_1_n) );
defparam Uadd_0_lut_l_2_n_1_n.IN_WIDTH = 26;
defparam Uadd_0_lut_l_2_n_1_n.PIPE_DEPTH = 1;

wire [27:0] tree_0_pp_l_3_n_0_n;
sadd_lpm Uadd_0_lut_l_3_n_0_n (.clk(clk), .ain(tree_0_pp_l_2_n_0_n), .bin(tree_0_pp_l_2_n_1_n), .res(tree_0_pp_l_3_n_0_n) );
defparam Uadd_0_lut_l_3_n_0_n.IN_WIDTH = 27;
defparam Uadd_0_lut_l_3_n_0_n.PIPE_DEPTH = 1;

wire [27:0] lut_val_0_n;
assign lut_val_0_n=tree_0_pp_l_3_n_0_n;


// ---- partial product adder tree ----

wire [23:0] lut_1_bit_0_fill;
wire [23:0] lut_1_bit_1_fill;
wire [23:0] lut_1_bit_2_fill;
wire [23:0] lut_1_bit_3_fill;
wire [23:0] lut_1_bit_4_fill;
wire [23:0] lut_1_bit_5_fill;
wire [23:0] lut_1_bit_6_fill;
wire [23:0] lut_1_bit_7_fill;
wire [23:0] lut_1_bit_8_fill;
wire [23:0] lut_1_bit_9_fill;
wire [23:0] lut_1_bit_10_fill;
wire [23:0] lut_1_bit_11_fill;
wire [23:0] lut_1_bit_12_fill;
wire [23:0] lut_1_bit_13_fill;
wire [23:0] lut_1_bit_14_fill;
wire [23:0] lut_1_bit_15_fill;
assign lut_1_bit_0_fill = {lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8], lut_val_1_n_0_pp[8],  lut_val_1_n_0_pp };
assign lut_1_bit_1_fill = {lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8], lut_val_1_n_1_pp[8],  lut_val_1_n_1_pp, 1'd0 };
assign lut_1_bit_2_fill = {lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8], lut_val_1_n_2_pp[8],  lut_val_1_n_2_pp, 2'd0 };
assign lut_1_bit_3_fill = {lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8], lut_val_1_n_3_pp[8],  lut_val_1_n_3_pp, 3'd0 };
assign lut_1_bit_4_fill = {lut_val_1_n_4_pp[8], lut_val_1_n_4_pp[8], lut_val_1_n_4_pp[8], lut_val_1_n_4_pp[8], lut_val_1_n_4_pp[8], lut_val_1_n_4_pp[8], lut_val_1_n_4_pp[8], lut_val_1_n_4_pp[8], lut_val_1_n_4_pp[8], lut_val_1_n_4_pp[8], lut_val_1_n_4_pp[8],  lut_val_1_n_4_pp, 4'd0 };
assign lut_1_bit_5_fill = {lut_val_1_n_5_pp[8], lut_val_1_n_5_pp[8], lut_val_1_n_5_pp[8], lut_val_1_n_5_pp[8], lut_val_1_n_5_pp[8], lut_val_1_n_5_pp[8], lut_val_1_n_5_pp[8], lut_val_1_n_5_pp[8], lut_val_1_n_5_pp[8], lut_val_1_n_5_pp[8],  lut_val_1_n_5_pp, 5'd0 };
assign lut_1_bit_6_fill = {lut_val_1_n_6_pp[8], lut_val_1_n_6_pp[8], lut_val_1_n_6_pp[8], lut_val_1_n_6_pp[8], lut_val_1_n_6_pp[8], lut_val_1_n_6_pp[8], lut_val_1_n_6_pp[8], lut_val_1_n_6_pp[8], lut_val_1_n_6_pp[8],  lut_val_1_n_6_pp, 6'd0 };
assign lut_1_bit_7_fill = {lut_val_1_n_7_pp[8], lut_val_1_n_7_pp[8], lut_val_1_n_7_pp[8], lut_val_1_n_7_pp[8], lut_val_1_n_7_pp[8], lut_val_1_n_7_pp[8], lut_val_1_n_7_pp[8], lut_val_1_n_7_pp[8],  lut_val_1_n_7_pp, 7'd0 };
assign lut_1_bit_8_fill = {lut_val_1_n_8_pp[8], lut_val_1_n_8_pp[8], lut_val_1_n_8_pp[8], lut_val_1_n_8_pp[8], lut_val_1_n_8_pp[8], lut_val_1_n_8_pp[8], lut_val_1_n_8_pp[8],  lut_val_1_n_8_pp, 8'd0 };
assign lut_1_bit_9_fill = {lut_val_1_n_9_pp[8], lut_val_1_n_9_pp[8], lut_val_1_n_9_pp[8], lut_val_1_n_9_pp[8], lut_val_1_n_9_pp[8], lut_val_1_n_9_pp[8],  lut_val_1_n_9_pp, 9'd0 };
assign lut_1_bit_10_fill = {lut_val_1_n_10_pp[8], lut_val_1_n_10_pp[8], lut_val_1_n_10_pp[8], lut_val_1_n_10_pp[8], lut_val_1_n_10_pp[8],  lut_val_1_n_10_pp, 10'd0 };
assign lut_1_bit_11_fill = {lut_val_1_n_11_pp[8], lut_val_1_n_11_pp[8], lut_val_1_n_11_pp[8], lut_val_1_n_11_pp[8],  lut_val_1_n_11_pp, 11'd0 };
assign lut_1_bit_12_fill = {lut_val_1_n_12_pp[8], lut_val_1_n_12_pp[8], lut_val_1_n_12_pp[8],  lut_val_1_n_12_pp, 12'd0 };
assign lut_1_bit_13_fill = {lut_val_1_n_13_pp[8], lut_val_1_n_13_pp[8],  lut_val_1_n_13_pp, 13'd0 };
assign lut_1_bit_14_fill = {lut_val_1_n_14_pp[8],  lut_val_1_n_14_pp, 14'd0 };
assign lut_1_bit_15_fill = { lut_val_1_n_15_pp, 15'd0 };
wire [24:0] tree_1_pp_l_0_n_0_n;
sadd_lpm Uadd_1_lut_l_0_n_0_n (.clk(clk), .ain(lut_1_bit_0_fill), .bin(lut_1_bit_1_fill), .res(tree_1_pp_l_0_n_0_n) );
defparam Uadd_1_lut_l_0_n_0_n.IN_WIDTH = 24;
defparam Uadd_1_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [24:0] tree_1_pp_l_0_n_1_n;
sadd_lpm Uadd_1_lut_l_0_n_1_n (.clk(clk), .ain(lut_1_bit_2_fill), .bin(lut_1_bit_3_fill), .res(tree_1_pp_l_0_n_1_n) );
defparam Uadd_1_lut_l_0_n_1_n.IN_WIDTH = 24;
defparam Uadd_1_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [24:0] tree_1_pp_l_0_n_2_n;
sadd_lpm Uadd_1_lut_l_0_n_2_n (.clk(clk), .ain(lut_1_bit_4_fill), .bin(lut_1_bit_5_fill), .res(tree_1_pp_l_0_n_2_n) );
defparam Uadd_1_lut_l_0_n_2_n.IN_WIDTH = 24;
defparam Uadd_1_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [24:0] tree_1_pp_l_0_n_3_n;
sadd_lpm Uadd_1_lut_l_0_n_3_n (.clk(clk), .ain(lut_1_bit_6_fill), .bin(lut_1_bit_7_fill), .res(tree_1_pp_l_0_n_3_n) );
defparam Uadd_1_lut_l_0_n_3_n.IN_WIDTH = 24;
defparam Uadd_1_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [24:0] tree_1_pp_l_0_n_4_n;
sadd_lpm Uadd_1_lut_l_0_n_4_n (.clk(clk), .ain(lut_1_bit_8_fill), .bin(lut_1_bit_9_fill), .res(tree_1_pp_l_0_n_4_n) );
defparam Uadd_1_lut_l_0_n_4_n.IN_WIDTH = 24;
defparam Uadd_1_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [24:0] tree_1_pp_l_0_n_5_n;
sadd_lpm Uadd_1_lut_l_0_n_5_n (.clk(clk), .ain(lut_1_bit_10_fill), .bin(lut_1_bit_11_fill), .res(tree_1_pp_l_0_n_5_n) );
defparam Uadd_1_lut_l_0_n_5_n.IN_WIDTH = 24;
defparam Uadd_1_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [24:0] tree_1_pp_l_0_n_6_n;
sadd_lpm Uadd_1_lut_l_0_n_6_n (.clk(clk), .ain(lut_1_bit_12_fill), .bin(lut_1_bit_13_fill), .res(tree_1_pp_l_0_n_6_n) );
defparam Uadd_1_lut_l_0_n_6_n.IN_WIDTH = 24;
defparam Uadd_1_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [24:0] tree_1_pp_l_0_n_7_n;
sadd_lpm Uadd_1_lut_l_0_n_7_n (.clk(clk), .ain(lut_1_bit_14_fill), .bin(lut_1_bit_15_fill), .res(tree_1_pp_l_0_n_7_n) );
defparam Uadd_1_lut_l_0_n_7_n.IN_WIDTH = 24;
defparam Uadd_1_lut_l_0_n_7_n.PIPE_DEPTH = 1;

wire [25:0] tree_1_pp_l_1_n_0_n;
sadd_lpm Uadd_1_lut_l_1_n_0_n (.clk(clk), .ain(tree_1_pp_l_0_n_0_n), .bin(tree_1_pp_l_0_n_1_n), .res(tree_1_pp_l_1_n_0_n) );
defparam Uadd_1_lut_l_1_n_0_n.IN_WIDTH = 25;
defparam Uadd_1_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [25:0] tree_1_pp_l_1_n_1_n;
sadd_lpm Uadd_1_lut_l_1_n_1_n (.clk(clk), .ain(tree_1_pp_l_0_n_2_n), .bin(tree_1_pp_l_0_n_3_n), .res(tree_1_pp_l_1_n_1_n) );
defparam Uadd_1_lut_l_1_n_1_n.IN_WIDTH = 25;
defparam Uadd_1_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [25:0] tree_1_pp_l_1_n_2_n;
sadd_lpm Uadd_1_lut_l_1_n_2_n (.clk(clk), .ain(tree_1_pp_l_0_n_4_n), .bin(tree_1_pp_l_0_n_5_n), .res(tree_1_pp_l_1_n_2_n) );
defparam Uadd_1_lut_l_1_n_2_n.IN_WIDTH = 25;
defparam Uadd_1_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [25:0] tree_1_pp_l_1_n_3_n;
sadd_lpm Uadd_1_lut_l_1_n_3_n (.clk(clk), .ain(tree_1_pp_l_0_n_6_n), .bin(tree_1_pp_l_0_n_7_n), .res(tree_1_pp_l_1_n_3_n) );
defparam Uadd_1_lut_l_1_n_3_n.IN_WIDTH = 25;
defparam Uadd_1_lut_l_1_n_3_n.PIPE_DEPTH = 1;

wire [26:0] tree_1_pp_l_2_n_0_n;
sadd_lpm Uadd_1_lut_l_2_n_0_n (.clk(clk), .ain(tree_1_pp_l_1_n_0_n), .bin(tree_1_pp_l_1_n_1_n), .res(tree_1_pp_l_2_n_0_n) );
defparam Uadd_1_lut_l_2_n_0_n.IN_WIDTH = 26;
defparam Uadd_1_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [26:0] tree_1_pp_l_2_n_1_n;
sadd_lpm Uadd_1_lut_l_2_n_1_n (.clk(clk), .ain(tree_1_pp_l_1_n_2_n), .bin(tree_1_pp_l_1_n_3_n), .res(tree_1_pp_l_2_n_1_n) );
defparam Uadd_1_lut_l_2_n_1_n.IN_WIDTH = 26;
defparam Uadd_1_lut_l_2_n_1_n.PIPE_DEPTH = 1;

wire [27:0] tree_1_pp_l_3_n_0_n;
sadd_lpm Uadd_1_lut_l_3_n_0_n (.clk(clk), .ain(tree_1_pp_l_2_n_0_n), .bin(tree_1_pp_l_2_n_1_n), .res(tree_1_pp_l_3_n_0_n) );
defparam Uadd_1_lut_l_3_n_0_n.IN_WIDTH = 27;
defparam Uadd_1_lut_l_3_n_0_n.PIPE_DEPTH = 1;

wire [27:0] lut_val_1_n;
assign lut_val_1_n=tree_1_pp_l_3_n_0_n;


// ---- final adder tree ----

wire [28:0] fin_atree_l_0_n_0_n;
sadd_lpm Uadd_l_0_n_0_n (.clk(clk), .ain(lut_val_0_n), .bin(lut_val_1_n), .res(fin_atree_l_0_n_0_n) );
defparam Uadd_l_0_n_0_n.IN_WIDTH = 28;
defparam Uadd_l_0_n_0_n.PIPE_DEPTH = 1;

wire [28:0] mac_res;
assign mac_res=fin_atree_l_0_n_0_n;
wire [28:0] atree_res;
mac_tl Umtl (.clk(clk), 
             .data_in(mac_res),
             .data_out(atree_res));
defparam Umtl.DATA_WIDTH = 29;

// ---- Adder Tree Complete ---- 
wire [28:0] fir_int_res;
assign fir_int_res = atree_res;

assign fir_result = fir_int_res[ACCUM_WIDTH-1:0];
endmodule
