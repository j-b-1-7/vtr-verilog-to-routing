`timescale 1ns / 1ns 
module system156(clk,resetn,boot_iaddr,boot_idata,boot_daddr,boot_ddata,reg_file_b_readdataout,processor_select);
	input clk;
	input resetn;
	input [8:0] processor_select;
	output [31:0] reg_file_b_readdataout;
	input [13:0] boot_iaddr;
	input [31:0] boot_idata;
	input [13:0] boot_daddr;
	input [31:0] boot_ddata;

	reg boot_iwe0;
	reg boot_dwe0;
	reg boot_iwe1;
	reg boot_dwe1;
	reg boot_iwe2;
	reg boot_dwe2;
	reg boot_iwe3;
	reg boot_dwe3;
	reg boot_iwe4;
	reg boot_dwe4;
	reg boot_iwe5;
	reg boot_dwe5;
	reg boot_iwe6;
	reg boot_dwe6;
	reg boot_iwe7;
	reg boot_dwe7;
	reg boot_iwe8;
	reg boot_dwe8;
	reg boot_iwe9;
	reg boot_dwe9;
	reg boot_iwe10;
	reg boot_dwe10;
	reg boot_iwe11;
	reg boot_dwe11;
	reg boot_iwe12;
	reg boot_dwe12;
	reg boot_iwe13;
	reg boot_dwe13;
	reg boot_iwe14;
	reg boot_dwe14;
	reg boot_iwe15;
	reg boot_dwe15;
	reg boot_iwe16;
	reg boot_dwe16;
	reg boot_iwe17;
	reg boot_dwe17;
	reg boot_iwe18;
	reg boot_dwe18;
	reg boot_iwe19;
	reg boot_dwe19;
	reg boot_iwe20;
	reg boot_dwe20;
	reg boot_iwe21;
	reg boot_dwe21;
	reg boot_iwe22;
	reg boot_dwe22;
	reg boot_iwe23;
	reg boot_dwe23;
	reg boot_iwe24;
	reg boot_dwe24;
	reg boot_iwe25;
	reg boot_dwe25;
	reg boot_iwe26;
	reg boot_dwe26;
	reg boot_iwe27;
	reg boot_dwe27;
	reg boot_iwe28;
	reg boot_dwe28;
	reg boot_iwe29;
	reg boot_dwe29;
	reg boot_iwe30;
	reg boot_dwe30;
	reg boot_iwe31;
	reg boot_dwe31;
	reg boot_iwe32;
	reg boot_dwe32;
	reg boot_iwe33;
	reg boot_dwe33;
	reg boot_iwe34;
	reg boot_dwe34;
	reg boot_iwe35;
	reg boot_dwe35;
	reg boot_iwe36;
	reg boot_dwe36;
	reg boot_iwe37;
	reg boot_dwe37;
	reg boot_iwe38;
	reg boot_dwe38;
	reg boot_iwe39;
	reg boot_dwe39;
	reg boot_iwe40;
	reg boot_dwe40;
	reg boot_iwe41;
	reg boot_dwe41;
	reg boot_iwe42;
	reg boot_dwe42;
	reg boot_iwe43;
	reg boot_dwe43;
	reg boot_iwe44;
	reg boot_dwe44;
	reg boot_iwe45;
	reg boot_dwe45;
	reg boot_iwe46;
	reg boot_dwe46;
	reg boot_iwe47;
	reg boot_dwe47;
	reg boot_iwe48;
	reg boot_dwe48;
	reg boot_iwe49;
	reg boot_dwe49;
	reg boot_iwe50;
	reg boot_dwe50;
	reg boot_iwe51;
	reg boot_dwe51;
	reg boot_iwe52;
	reg boot_dwe52;
	reg boot_iwe53;
	reg boot_dwe53;
	reg boot_iwe54;
	reg boot_dwe54;
	reg boot_iwe55;
	reg boot_dwe55;
	reg boot_iwe56;
	reg boot_dwe56;
	reg boot_iwe57;
	reg boot_dwe57;
	reg boot_iwe58;
	reg boot_dwe58;
	reg boot_iwe59;
	reg boot_dwe59;
	reg boot_iwe60;
	reg boot_dwe60;
	reg boot_iwe61;
	reg boot_dwe61;
	reg boot_iwe62;
	reg boot_dwe62;
	reg boot_iwe63;
	reg boot_dwe63;
	reg boot_iwe64;
	reg boot_dwe64;
	reg boot_iwe65;
	reg boot_dwe65;
	reg boot_iwe66;
	reg boot_dwe66;
	reg boot_iwe67;
	reg boot_dwe67;
	reg boot_iwe68;
	reg boot_dwe68;
	reg boot_iwe69;
	reg boot_dwe69;
	reg boot_iwe70;
	reg boot_dwe70;
	reg boot_iwe71;
	reg boot_dwe71;
	reg boot_iwe72;
	reg boot_dwe72;
	reg boot_iwe73;
	reg boot_dwe73;
	reg boot_iwe74;
	reg boot_dwe74;
	reg boot_iwe75;
	reg boot_dwe75;
	reg boot_iwe76;
	reg boot_dwe76;
	reg boot_iwe77;
	reg boot_dwe77;
	reg boot_iwe78;
	reg boot_dwe78;
	reg boot_iwe79;
	reg boot_dwe79;
	reg boot_iwe80;
	reg boot_dwe80;
	reg boot_iwe81;
	reg boot_dwe81;
	reg boot_iwe82;
	reg boot_dwe82;
	reg boot_iwe83;
	reg boot_dwe83;
	reg boot_iwe84;
	reg boot_dwe84;
	reg boot_iwe85;
	reg boot_dwe85;
	reg boot_iwe86;
	reg boot_dwe86;
	reg boot_iwe87;
	reg boot_dwe87;
	reg boot_iwe88;
	reg boot_dwe88;
	reg boot_iwe89;
	reg boot_dwe89;
	reg boot_iwe90;
	reg boot_dwe90;
	reg boot_iwe91;
	reg boot_dwe91;
	reg boot_iwe92;
	reg boot_dwe92;
	reg boot_iwe93;
	reg boot_dwe93;
	reg boot_iwe94;
	reg boot_dwe94;
	reg boot_iwe95;
	reg boot_dwe95;
	reg boot_iwe96;
	reg boot_dwe96;
	reg boot_iwe97;
	reg boot_dwe97;
	reg boot_iwe98;
	reg boot_dwe98;
	reg boot_iwe99;
	reg boot_dwe99;
	reg boot_iwe100;
	reg boot_dwe100;
	reg boot_iwe101;
	reg boot_dwe101;
	reg boot_iwe102;
	reg boot_dwe102;
	reg boot_iwe103;
	reg boot_dwe103;
	reg boot_iwe104;
	reg boot_dwe104;
	reg boot_iwe105;
	reg boot_dwe105;
	reg boot_iwe106;
	reg boot_dwe106;
	reg boot_iwe107;
	reg boot_dwe107;
	reg boot_iwe108;
	reg boot_dwe108;
	reg boot_iwe109;
	reg boot_dwe109;
	reg boot_iwe110;
	reg boot_dwe110;
	reg boot_iwe111;
	reg boot_dwe111;
	reg boot_iwe112;
	reg boot_dwe112;
	reg boot_iwe113;
	reg boot_dwe113;
	reg boot_iwe114;
	reg boot_dwe114;
	reg boot_iwe115;
	reg boot_dwe115;
	reg boot_iwe116;
	reg boot_dwe116;
	reg boot_iwe117;
	reg boot_dwe117;
	reg boot_iwe118;
	reg boot_dwe118;
	reg boot_iwe119;
	reg boot_dwe119;
	reg boot_iwe120;
	reg boot_dwe120;
	reg boot_iwe121;
	reg boot_dwe121;
	reg boot_iwe122;
	reg boot_dwe122;
	reg boot_iwe123;
	reg boot_dwe123;
	reg boot_iwe124;
	reg boot_dwe124;
	reg boot_iwe125;
	reg boot_dwe125;
	reg boot_iwe126;
	reg boot_dwe126;
	reg boot_iwe127;
	reg boot_dwe127;
	reg boot_iwe128;
	reg boot_dwe128;
	reg boot_iwe129;
	reg boot_dwe129;
	reg boot_iwe130;
	reg boot_dwe130;
	reg boot_iwe131;
	reg boot_dwe131;
	reg boot_iwe132;
	reg boot_dwe132;
	reg boot_iwe133;
	reg boot_dwe133;
	reg boot_iwe134;
	reg boot_dwe134;
	reg boot_iwe135;
	reg boot_dwe135;
	reg boot_iwe136;
	reg boot_dwe136;
	reg boot_iwe137;
	reg boot_dwe137;
	reg boot_iwe138;
	reg boot_dwe138;
	reg boot_iwe139;
	reg boot_dwe139;
	reg boot_iwe140;
	reg boot_dwe140;
	reg boot_iwe141;
	reg boot_dwe141;
	reg boot_iwe142;
	reg boot_dwe142;
	reg boot_iwe143;
	reg boot_dwe143;
	reg boot_iwe144;
	reg boot_dwe144;
	reg boot_iwe145;
	reg boot_dwe145;
	reg boot_iwe146;
	reg boot_dwe146;
	reg boot_iwe147;
	reg boot_dwe147;
	reg boot_iwe148;
	reg boot_dwe148;
	reg boot_iwe149;
	reg boot_dwe149;
	reg boot_iwe150;
	reg boot_dwe150;
	reg boot_iwe151;
	reg boot_dwe151;
	reg boot_iwe152;
	reg boot_dwe152;
	reg boot_iwe153;
	reg boot_dwe153;
	reg boot_iwe154;
	reg boot_dwe154;
	reg boot_iwe155;
	reg boot_dwe155;
 
	 //Processor 0 control and data signals
	wire rdProc0South;
	wire emptyProc0South;
	wire [31:0] dataInProc0South;

	 //Processor 0 control and data signals
	wire wrProc0South;
	wire fullProc0South;
	wire [31:0] dataOutProc0South;
	
	//Processor 0 control and data signals
	wire rdProc0East;
	wire emptyProc0East;
	wire [31:0] dataInProc0East;

	 //Processor 0 control and data signals
	wire wrProc0East;
	wire fullProc0East;
	wire [31:0] dataOutProc0East;
	
	 //Processor 1 control and data signals
	wire rdProc1South;
	wire emptyProc1South;
	wire [31:0] dataInProc1South;

	 //Processor 1 control and data signals
	wire wrProc1South;
	wire fullProc1South;
	wire [31:0] dataOutProc1South;

	 //Processor 1 control and data signals
	wire rdProc1East;
	wire emptyProc1East;
	wire [31:0] dataInProc1East;
	
	//Processor 1 control and data signals
	wire wrProc1East;
	wire fullProc1East;
	wire [31:0] dataOutProc1East;

	 //Processor 1 control and data signals
	wire rdProc1West;
	wire emptyProc1West;
	wire [31:0] dataInProc1West;
	
	//Processor 1 control and data signals
	wire wrProc1West;
	wire fullProc1West;
	wire [31:0] dataOutProc1West;
	
	 //Processor 2 control and data signals
	wire rdProc2South;
	wire emptyProc2South;
	wire [31:0] dataInProc2South;

	 //Processor 2 control and data signals
	wire wrProc2South;
	wire fullProc2South;
	wire [31:0] dataOutProc2South;

	 //Processor 2 control and data signals
	wire rdProc2East;
	wire emptyProc2East;
	wire [31:0] dataInProc2East;
	
	//Processor 2 control and data signals
	wire wrProc2East;
	wire fullProc2East;
	wire [31:0] dataOutProc2East;

	 //Processor 2 control and data signals
	wire rdProc2West;
	wire emptyProc2West;
	wire [31:0] dataInProc2West;
	
	//Processor 2 control and data signals
	wire wrProc2West;
	wire fullProc2West;
	wire [31:0] dataOutProc2West;
	
	 //Processor 3 control and data signals
	wire rdProc3South;
	wire emptyProc3South;
	wire [31:0] dataInProc3South;

	 //Processor 3 control and data signals
	wire wrProc3South;
	wire fullProc3South;
	wire [31:0] dataOutProc3South;

	 //Processor 3 control and data signals
	wire rdProc3East;
	wire emptyProc3East;
	wire [31:0] dataInProc3East;
	
	//Processor 3 control and data signals
	wire wrProc3East;
	wire fullProc3East;
	wire [31:0] dataOutProc3East;

	 //Processor 3 control and data signals
	wire rdProc3West;
	wire emptyProc3West;
	wire [31:0] dataInProc3West;
	
	//Processor 3 control and data signals
	wire wrProc3West;
	wire fullProc3West;
	wire [31:0] dataOutProc3West;
	
	 //Processor 4 control and data signals
	wire rdProc4South;
	wire emptyProc4South;
	wire [31:0] dataInProc4South;

	 //Processor 4 control and data signals
	wire wrProc4South;
	wire fullProc4South;
	wire [31:0] dataOutProc4South;

	 //Processor 4 control and data signals
	wire rdProc4East;
	wire emptyProc4East;
	wire [31:0] dataInProc4East;
	
	//Processor 4 control and data signals
	wire wrProc4East;
	wire fullProc4East;
	wire [31:0] dataOutProc4East;

	 //Processor 4 control and data signals
	wire rdProc4West;
	wire emptyProc4West;
	wire [31:0] dataInProc4West;
	
	//Processor 4 control and data signals
	wire wrProc4West;
	wire fullProc4West;
	wire [31:0] dataOutProc4West;
	
	 //Processor 5 control and data signals
	wire rdProc5South;
	wire emptyProc5South;
	wire [31:0] dataInProc5South;

	 //Processor 5 control and data signals
	wire wrProc5South;
	wire fullProc5South;
	wire [31:0] dataOutProc5South;

	 //Processor 5 control and data signals
	wire rdProc5East;
	wire emptyProc5East;
	wire [31:0] dataInProc5East;
	
	//Processor 5 control and data signals
	wire wrProc5East;
	wire fullProc5East;
	wire [31:0] dataOutProc5East;

	 //Processor 5 control and data signals
	wire rdProc5West;
	wire emptyProc5West;
	wire [31:0] dataInProc5West;
	
	//Processor 5 control and data signals
	wire wrProc5West;
	wire fullProc5West;
	wire [31:0] dataOutProc5West;
	
	 //Processor 6 control and data signals
	wire rdProc6South;
	wire emptyProc6South;
	wire [31:0] dataInProc6South;

	 //Processor 6 control and data signals
	wire wrProc6South;
	wire fullProc6South;
	wire [31:0] dataOutProc6South;

	 //Processor 6 control and data signals
	wire rdProc6East;
	wire emptyProc6East;
	wire [31:0] dataInProc6East;
	
	//Processor 6 control and data signals
	wire wrProc6East;
	wire fullProc6East;
	wire [31:0] dataOutProc6East;

	 //Processor 6 control and data signals
	wire rdProc6West;
	wire emptyProc6West;
	wire [31:0] dataInProc6West;
	
	//Processor 6 control and data signals
	wire wrProc6West;
	wire fullProc6West;
	wire [31:0] dataOutProc6West;
	
	 //Processor 7 control and data signals
	wire rdProc7South;
	wire emptyProc7South;
	wire [31:0] dataInProc7South;

	 //Processor 7 control and data signals
	wire wrProc7South;
	wire fullProc7South;
	wire [31:0] dataOutProc7South;

	 //Processor 7 control and data signals
	wire rdProc7East;
	wire emptyProc7East;
	wire [31:0] dataInProc7East;
	
	//Processor 7 control and data signals
	wire wrProc7East;
	wire fullProc7East;
	wire [31:0] dataOutProc7East;

	 //Processor 7 control and data signals
	wire rdProc7West;
	wire emptyProc7West;
	wire [31:0] dataInProc7West;
	
	//Processor 7 control and data signals
	wire wrProc7West;
	wire fullProc7West;
	wire [31:0] dataOutProc7West;
	
	 //Processor 8 control and data signals
	wire rdProc8South;
	wire emptyProc8South;
	wire [31:0] dataInProc8South;

	 //Processor 8 control and data signals
	wire wrProc8South;
	wire fullProc8South;
	wire [31:0] dataOutProc8South;

	 //Processor 8 control and data signals
	wire rdProc8East;
	wire emptyProc8East;
	wire [31:0] dataInProc8East;
	
	//Processor 8 control and data signals
	wire wrProc8East;
	wire fullProc8East;
	wire [31:0] dataOutProc8East;

	 //Processor 8 control and data signals
	wire rdProc8West;
	wire emptyProc8West;
	wire [31:0] dataInProc8West;
	
	//Processor 8 control and data signals
	wire wrProc8West;
	wire fullProc8West;
	wire [31:0] dataOutProc8West;
	
	 //Processor 9 control and data signals
	wire rdProc9South;
	wire emptyProc9South;
	wire [31:0] dataInProc9South;

	 //Processor 9 control and data signals
	wire wrProc9South;
	wire fullProc9South;
	wire [31:0] dataOutProc9South;

	 //Processor 9 control and data signals
	wire rdProc9East;
	wire emptyProc9East;
	wire [31:0] dataInProc9East;
	
	//Processor 9 control and data signals
	wire wrProc9East;
	wire fullProc9East;
	wire [31:0] dataOutProc9East;

	 //Processor 9 control and data signals
	wire rdProc9West;
	wire emptyProc9West;
	wire [31:0] dataInProc9West;
	
	//Processor 9 control and data signals
	wire wrProc9West;
	wire fullProc9West;
	wire [31:0] dataOutProc9West;
	
	 //Processor 10 control and data signals
	wire rdProc10South;
	wire emptyProc10South;
	wire [31:0] dataInProc10South;

	 //Processor 10 control and data signals
	wire wrProc10South;
	wire fullProc10South;
	wire [31:0] dataOutProc10South;

	 //Processor 10 control and data signals
	wire rdProc10East;
	wire emptyProc10East;
	wire [31:0] dataInProc10East;
	
	//Processor 10 control and data signals
	wire wrProc10East;
	wire fullProc10East;
	wire [31:0] dataOutProc10East;

	 //Processor 10 control and data signals
	wire rdProc10West;
	wire emptyProc10West;
	wire [31:0] dataInProc10West;
	
	//Processor 10 control and data signals
	wire wrProc10West;
	wire fullProc10West;
	wire [31:0] dataOutProc10West;
	
	 //Processor 11 control and data signals
	wire rdProc11South;
	wire emptyProc11South;
	wire [31:0] dataInProc11South;

	 //Processor 11 control and data signals
	wire wrProc11South;
	wire fullProc11South;
	wire [31:0] dataOutProc11South;

	 //Processor 11 control and data signals
	wire rdProc11East;
	wire emptyProc11East;
	wire [31:0] dataInProc11East;
	
	//Processor 11 control and data signals
	wire wrProc11East;
	wire fullProc11East;
	wire [31:0] dataOutProc11East;

	 //Processor 11 control and data signals
	wire rdProc11West;
	wire emptyProc11West;
	wire [31:0] dataInProc11West;
	
	//Processor 11 control and data signals
	wire wrProc11West;
	wire fullProc11West;
	wire [31:0] dataOutProc11West;
	
	 //Processor 12 control and data signals
	wire rdProc12South;
	wire emptyProc12South;
	wire [31:0] dataInProc12South;

	 //Processor 12 control and data signals
	wire wrProc12South;
	wire fullProc12South;
	wire [31:0] dataOutProc12South;
	
	 //Processor 12 control and data signals
	wire wrProc12West;
	wire fullProc12West;
	wire [31:0] dataOutProc12West;

	 //Processor 12 control and data signals
	wire rdProc12West;
	wire emptyProc12West;
	wire [31:0] dataInProc12West;

	//Processor 13 control and data signals
	wire wrProc13North;
	wire fullProc13North;
	wire [31:0] dataOutProc13North;

	 //Processor 13 control and data signals
	wire rdProc13North;
	wire emptyProc13North;
	wire [31:0] dataInProc13North;
	
	 //Processor 13 control and data signals
	wire rdProc13South;
	wire emptyProc13South;
	wire [31:0] dataInProc13South;
	
	 //Processor 13 control and data signals
	wire wrProc13South;
	wire fullProc13South;
	wire [31:0] dataOutProc13South;
	
	 //Processor 13 control and data signals
	wire rdProc13East;
	wire emptyProc13East;
	wire [31:0] dataInProc13East;

	 //Processor 13 control and data signals
	wire wrProc13East;
	wire fullProc13East;
	wire [31:0] dataOutProc13East;

	//Processor 14 control and data signals
	wire rdProc14North;
	wire emptyProc14North;
	wire [31:0] dataInProc14North;

	 //Processor 14 control and data signals
	wire wrProc14North;
	wire fullProc14North;
	wire [31:0] dataOutProc14North;

	 //Processor 14 control and data signals
	wire rdProc14South;
	wire emptyProc14South;
	wire [31:0] dataInProc14South;
	
	 //Processor 14 control and data signals
	wire wrProc14South;
	wire fullProc14South;
	wire [31:0] dataOutProc14South;

	 //Processor 14 control and data signals
	wire rdProc14East;
	wire emptyProc14East;
	wire [31:0] dataInProc14East;
	
	 //Processor 14 control and data signals
	wire wrProc14East;
	wire fullProc14East;
	wire [31:0] dataOutProc14East;

	 //Processor 14 control and data signals
	wire rdProc14West;
	wire emptyProc14West;
	wire [31:0] dataInProc14West;

	 //Processor 14 control and data signals
	wire wrProc14West;
	wire fullProc14West;
	wire [31:0] dataOutProc14West;

	//Processor 15 control and data signals
	wire rdProc15North;
	wire emptyProc15North;
	wire [31:0] dataInProc15North;

	 //Processor 15 control and data signals
	wire wrProc15North;
	wire fullProc15North;
	wire [31:0] dataOutProc15North;

	 //Processor 15 control and data signals
	wire rdProc15South;
	wire emptyProc15South;
	wire [31:0] dataInProc15South;
	
	 //Processor 15 control and data signals
	wire wrProc15South;
	wire fullProc15South;
	wire [31:0] dataOutProc15South;

	 //Processor 15 control and data signals
	wire rdProc15East;
	wire emptyProc15East;
	wire [31:0] dataInProc15East;
	
	 //Processor 15 control and data signals
	wire wrProc15East;
	wire fullProc15East;
	wire [31:0] dataOutProc15East;

	 //Processor 15 control and data signals
	wire rdProc15West;
	wire emptyProc15West;
	wire [31:0] dataInProc15West;

	 //Processor 15 control and data signals
	wire wrProc15West;
	wire fullProc15West;
	wire [31:0] dataOutProc15West;

	//Processor 16 control and data signals
	wire rdProc16North;
	wire emptyProc16North;
	wire [31:0] dataInProc16North;

	 //Processor 16 control and data signals
	wire wrProc16North;
	wire fullProc16North;
	wire [31:0] dataOutProc16North;

	 //Processor 16 control and data signals
	wire rdProc16South;
	wire emptyProc16South;
	wire [31:0] dataInProc16South;
	
	 //Processor 16 control and data signals
	wire wrProc16South;
	wire fullProc16South;
	wire [31:0] dataOutProc16South;

	 //Processor 16 control and data signals
	wire rdProc16East;
	wire emptyProc16East;
	wire [31:0] dataInProc16East;
	
	 //Processor 16 control and data signals
	wire wrProc16East;
	wire fullProc16East;
	wire [31:0] dataOutProc16East;

	 //Processor 16 control and data signals
	wire rdProc16West;
	wire emptyProc16West;
	wire [31:0] dataInProc16West;

	 //Processor 16 control and data signals
	wire wrProc16West;
	wire fullProc16West;
	wire [31:0] dataOutProc16West;

	//Processor 17 control and data signals
	wire rdProc17North;
	wire emptyProc17North;
	wire [31:0] dataInProc17North;

	 //Processor 17 control and data signals
	wire wrProc17North;
	wire fullProc17North;
	wire [31:0] dataOutProc17North;

	 //Processor 17 control and data signals
	wire rdProc17South;
	wire emptyProc17South;
	wire [31:0] dataInProc17South;
	
	 //Processor 17 control and data signals
	wire wrProc17South;
	wire fullProc17South;
	wire [31:0] dataOutProc17South;

	 //Processor 17 control and data signals
	wire rdProc17East;
	wire emptyProc17East;
	wire [31:0] dataInProc17East;
	
	 //Processor 17 control and data signals
	wire wrProc17East;
	wire fullProc17East;
	wire [31:0] dataOutProc17East;

	 //Processor 17 control and data signals
	wire rdProc17West;
	wire emptyProc17West;
	wire [31:0] dataInProc17West;

	 //Processor 17 control and data signals
	wire wrProc17West;
	wire fullProc17West;
	wire [31:0] dataOutProc17West;

	//Processor 18 control and data signals
	wire rdProc18North;
	wire emptyProc18North;
	wire [31:0] dataInProc18North;

	 //Processor 18 control and data signals
	wire wrProc18North;
	wire fullProc18North;
	wire [31:0] dataOutProc18North;

	 //Processor 18 control and data signals
	wire rdProc18South;
	wire emptyProc18South;
	wire [31:0] dataInProc18South;
	
	 //Processor 18 control and data signals
	wire wrProc18South;
	wire fullProc18South;
	wire [31:0] dataOutProc18South;

	 //Processor 18 control and data signals
	wire rdProc18East;
	wire emptyProc18East;
	wire [31:0] dataInProc18East;
	
	 //Processor 18 control and data signals
	wire wrProc18East;
	wire fullProc18East;
	wire [31:0] dataOutProc18East;

	 //Processor 18 control and data signals
	wire rdProc18West;
	wire emptyProc18West;
	wire [31:0] dataInProc18West;

	 //Processor 18 control and data signals
	wire wrProc18West;
	wire fullProc18West;
	wire [31:0] dataOutProc18West;

	//Processor 19 control and data signals
	wire rdProc19North;
	wire emptyProc19North;
	wire [31:0] dataInProc19North;

	 //Processor 19 control and data signals
	wire wrProc19North;
	wire fullProc19North;
	wire [31:0] dataOutProc19North;

	 //Processor 19 control and data signals
	wire rdProc19South;
	wire emptyProc19South;
	wire [31:0] dataInProc19South;
	
	 //Processor 19 control and data signals
	wire wrProc19South;
	wire fullProc19South;
	wire [31:0] dataOutProc19South;

	 //Processor 19 control and data signals
	wire rdProc19East;
	wire emptyProc19East;
	wire [31:0] dataInProc19East;
	
	 //Processor 19 control and data signals
	wire wrProc19East;
	wire fullProc19East;
	wire [31:0] dataOutProc19East;

	 //Processor 19 control and data signals
	wire rdProc19West;
	wire emptyProc19West;
	wire [31:0] dataInProc19West;

	 //Processor 19 control and data signals
	wire wrProc19West;
	wire fullProc19West;
	wire [31:0] dataOutProc19West;

	//Processor 20 control and data signals
	wire rdProc20North;
	wire emptyProc20North;
	wire [31:0] dataInProc20North;

	 //Processor 20 control and data signals
	wire wrProc20North;
	wire fullProc20North;
	wire [31:0] dataOutProc20North;

	 //Processor 20 control and data signals
	wire rdProc20South;
	wire emptyProc20South;
	wire [31:0] dataInProc20South;
	
	 //Processor 20 control and data signals
	wire wrProc20South;
	wire fullProc20South;
	wire [31:0] dataOutProc20South;

	 //Processor 20 control and data signals
	wire rdProc20East;
	wire emptyProc20East;
	wire [31:0] dataInProc20East;
	
	 //Processor 20 control and data signals
	wire wrProc20East;
	wire fullProc20East;
	wire [31:0] dataOutProc20East;

	 //Processor 20 control and data signals
	wire rdProc20West;
	wire emptyProc20West;
	wire [31:0] dataInProc20West;

	 //Processor 20 control and data signals
	wire wrProc20West;
	wire fullProc20West;
	wire [31:0] dataOutProc20West;

	//Processor 21 control and data signals
	wire rdProc21North;
	wire emptyProc21North;
	wire [31:0] dataInProc21North;

	 //Processor 21 control and data signals
	wire wrProc21North;
	wire fullProc21North;
	wire [31:0] dataOutProc21North;

	 //Processor 21 control and data signals
	wire rdProc21South;
	wire emptyProc21South;
	wire [31:0] dataInProc21South;
	
	 //Processor 21 control and data signals
	wire wrProc21South;
	wire fullProc21South;
	wire [31:0] dataOutProc21South;

	 //Processor 21 control and data signals
	wire rdProc21East;
	wire emptyProc21East;
	wire [31:0] dataInProc21East;
	
	 //Processor 21 control and data signals
	wire wrProc21East;
	wire fullProc21East;
	wire [31:0] dataOutProc21East;

	 //Processor 21 control and data signals
	wire rdProc21West;
	wire emptyProc21West;
	wire [31:0] dataInProc21West;

	 //Processor 21 control and data signals
	wire wrProc21West;
	wire fullProc21West;
	wire [31:0] dataOutProc21West;

	//Processor 22 control and data signals
	wire rdProc22North;
	wire emptyProc22North;
	wire [31:0] dataInProc22North;

	 //Processor 22 control and data signals
	wire wrProc22North;
	wire fullProc22North;
	wire [31:0] dataOutProc22North;

	 //Processor 22 control and data signals
	wire rdProc22South;
	wire emptyProc22South;
	wire [31:0] dataInProc22South;
	
	 //Processor 22 control and data signals
	wire wrProc22South;
	wire fullProc22South;
	wire [31:0] dataOutProc22South;

	 //Processor 22 control and data signals
	wire rdProc22East;
	wire emptyProc22East;
	wire [31:0] dataInProc22East;
	
	 //Processor 22 control and data signals
	wire wrProc22East;
	wire fullProc22East;
	wire [31:0] dataOutProc22East;

	 //Processor 22 control and data signals
	wire rdProc22West;
	wire emptyProc22West;
	wire [31:0] dataInProc22West;

	 //Processor 22 control and data signals
	wire wrProc22West;
	wire fullProc22West;
	wire [31:0] dataOutProc22West;

	//Processor 23 control and data signals
	wire rdProc23North;
	wire emptyProc23North;
	wire [31:0] dataInProc23North;

	 //Processor 23 control and data signals
	wire wrProc23North;
	wire fullProc23North;
	wire [31:0] dataOutProc23North;

	 //Processor 23 control and data signals
	wire rdProc23South;
	wire emptyProc23South;
	wire [31:0] dataInProc23South;
	
	 //Processor 23 control and data signals
	wire wrProc23South;
	wire fullProc23South;
	wire [31:0] dataOutProc23South;

	 //Processor 23 control and data signals
	wire rdProc23East;
	wire emptyProc23East;
	wire [31:0] dataInProc23East;
	
	 //Processor 23 control and data signals
	wire wrProc23East;
	wire fullProc23East;
	wire [31:0] dataOutProc23East;

	 //Processor 23 control and data signals
	wire rdProc23West;
	wire emptyProc23West;
	wire [31:0] dataInProc23West;

	 //Processor 23 control and data signals
	wire wrProc23West;
	wire fullProc23West;
	wire [31:0] dataOutProc23West;

	//Processor 24 control and data signals
	wire rdProc24North;
	wire emptyProc24North;
	wire [31:0] dataInProc24North;

	 //Processor 24 control and data signals
	wire wrProc24North;
	wire fullProc24North;
	wire [31:0] dataOutProc24North;

	 //Processor 24 control and data signals
	wire rdProc24South;
	wire emptyProc24South;
	wire [31:0] dataInProc24South;
	
	 //Processor 24 control and data signals
	wire wrProc24South;
	wire fullProc24South;
	wire [31:0] dataOutProc24South;

	 //Processor 24 control and data signals
	wire rdProc24East;
	wire emptyProc24East;
	wire [31:0] dataInProc24East;
	
	 //Processor 24 control and data signals
	wire wrProc24East;
	wire fullProc24East;
	wire [31:0] dataOutProc24East;

	 //Processor 24 control and data signals
	wire rdProc24West;
	wire emptyProc24West;
	wire [31:0] dataInProc24West;

	 //Processor 24 control and data signals
	wire wrProc24West;
	wire fullProc24West;
	wire [31:0] dataOutProc24West;

	//Processor 25 control and data signals
	wire wrProc25North;
	wire fullProc25North;
	wire [31:0] dataOutProc25North;

	//Processor 25 control and data signals
        wire rdProc25North;
        wire emptyProc25North;
        wire [31:0] dataInProc25North;

	//Processor 25 control and data signals
	wire rdProc25South;
	wire emptyProc25South;
	wire [31:0] dataInProc25South;
		
	 //Processor 25 control and data signals
	wire wrProc25South;
	wire fullProc25South;
	wire [31:0] dataOutProc25South;

	 //Processor 25 control and data signals
	wire wrProc25West;
	wire fullProc25West;
	wire [31:0] dataOutProc25West;
	
	 //Processor 25 control and data signals
	wire rdProc25West;
	wire emptyProc25West;
	wire [31:0] dataInProc25West;

	//Processor 26 control and data signals
	wire wrProc26North;
	wire fullProc26North;
	wire [31:0] dataOutProc26North;

	 //Processor 26 control and data signals
	wire rdProc26North;
	wire emptyProc26North;
	wire [31:0] dataInProc26North;
	
	 //Processor 26 control and data signals
	wire rdProc26South;
	wire emptyProc26South;
	wire [31:0] dataInProc26South;
	
	 //Processor 26 control and data signals
	wire wrProc26South;
	wire fullProc26South;
	wire [31:0] dataOutProc26South;
	
	 //Processor 26 control and data signals
	wire rdProc26East;
	wire emptyProc26East;
	wire [31:0] dataInProc26East;

	 //Processor 26 control and data signals
	wire wrProc26East;
	wire fullProc26East;
	wire [31:0] dataOutProc26East;

	//Processor 27 control and data signals
	wire rdProc27North;
	wire emptyProc27North;
	wire [31:0] dataInProc27North;

	 //Processor 27 control and data signals
	wire wrProc27North;
	wire fullProc27North;
	wire [31:0] dataOutProc27North;

	 //Processor 27 control and data signals
	wire rdProc27South;
	wire emptyProc27South;
	wire [31:0] dataInProc27South;
	
	 //Processor 27 control and data signals
	wire wrProc27South;
	wire fullProc27South;
	wire [31:0] dataOutProc27South;

	 //Processor 27 control and data signals
	wire rdProc27East;
	wire emptyProc27East;
	wire [31:0] dataInProc27East;
	
	 //Processor 27 control and data signals
	wire wrProc27East;
	wire fullProc27East;
	wire [31:0] dataOutProc27East;

	 //Processor 27 control and data signals
	wire rdProc27West;
	wire emptyProc27West;
	wire [31:0] dataInProc27West;

	 //Processor 27 control and data signals
	wire wrProc27West;
	wire fullProc27West;
	wire [31:0] dataOutProc27West;

	//Processor 28 control and data signals
	wire rdProc28North;
	wire emptyProc28North;
	wire [31:0] dataInProc28North;

	 //Processor 28 control and data signals
	wire wrProc28North;
	wire fullProc28North;
	wire [31:0] dataOutProc28North;

	 //Processor 28 control and data signals
	wire rdProc28South;
	wire emptyProc28South;
	wire [31:0] dataInProc28South;
	
	 //Processor 28 control and data signals
	wire wrProc28South;
	wire fullProc28South;
	wire [31:0] dataOutProc28South;

	 //Processor 28 control and data signals
	wire rdProc28East;
	wire emptyProc28East;
	wire [31:0] dataInProc28East;
	
	 //Processor 28 control and data signals
	wire wrProc28East;
	wire fullProc28East;
	wire [31:0] dataOutProc28East;

	 //Processor 28 control and data signals
	wire rdProc28West;
	wire emptyProc28West;
	wire [31:0] dataInProc28West;

	 //Processor 28 control and data signals
	wire wrProc28West;
	wire fullProc28West;
	wire [31:0] dataOutProc28West;

	//Processor 29 control and data signals
	wire rdProc29North;
	wire emptyProc29North;
	wire [31:0] dataInProc29North;

	 //Processor 29 control and data signals
	wire wrProc29North;
	wire fullProc29North;
	wire [31:0] dataOutProc29North;

	 //Processor 29 control and data signals
	wire rdProc29South;
	wire emptyProc29South;
	wire [31:0] dataInProc29South;
	
	 //Processor 29 control and data signals
	wire wrProc29South;
	wire fullProc29South;
	wire [31:0] dataOutProc29South;

	 //Processor 29 control and data signals
	wire rdProc29East;
	wire emptyProc29East;
	wire [31:0] dataInProc29East;
	
	 //Processor 29 control and data signals
	wire wrProc29East;
	wire fullProc29East;
	wire [31:0] dataOutProc29East;

	 //Processor 29 control and data signals
	wire rdProc29West;
	wire emptyProc29West;
	wire [31:0] dataInProc29West;

	 //Processor 29 control and data signals
	wire wrProc29West;
	wire fullProc29West;
	wire [31:0] dataOutProc29West;

	//Processor 30 control and data signals
	wire rdProc30North;
	wire emptyProc30North;
	wire [31:0] dataInProc30North;

	 //Processor 30 control and data signals
	wire wrProc30North;
	wire fullProc30North;
	wire [31:0] dataOutProc30North;

	 //Processor 30 control and data signals
	wire rdProc30South;
	wire emptyProc30South;
	wire [31:0] dataInProc30South;
	
	 //Processor 30 control and data signals
	wire wrProc30South;
	wire fullProc30South;
	wire [31:0] dataOutProc30South;

	 //Processor 30 control and data signals
	wire rdProc30East;
	wire emptyProc30East;
	wire [31:0] dataInProc30East;
	
	 //Processor 30 control and data signals
	wire wrProc30East;
	wire fullProc30East;
	wire [31:0] dataOutProc30East;

	 //Processor 30 control and data signals
	wire rdProc30West;
	wire emptyProc30West;
	wire [31:0] dataInProc30West;

	 //Processor 30 control and data signals
	wire wrProc30West;
	wire fullProc30West;
	wire [31:0] dataOutProc30West;

	//Processor 31 control and data signals
	wire rdProc31North;
	wire emptyProc31North;
	wire [31:0] dataInProc31North;

	 //Processor 31 control and data signals
	wire wrProc31North;
	wire fullProc31North;
	wire [31:0] dataOutProc31North;

	 //Processor 31 control and data signals
	wire rdProc31South;
	wire emptyProc31South;
	wire [31:0] dataInProc31South;
	
	 //Processor 31 control and data signals
	wire wrProc31South;
	wire fullProc31South;
	wire [31:0] dataOutProc31South;

	 //Processor 31 control and data signals
	wire rdProc31East;
	wire emptyProc31East;
	wire [31:0] dataInProc31East;
	
	 //Processor 31 control and data signals
	wire wrProc31East;
	wire fullProc31East;
	wire [31:0] dataOutProc31East;

	 //Processor 31 control and data signals
	wire rdProc31West;
	wire emptyProc31West;
	wire [31:0] dataInProc31West;

	 //Processor 31 control and data signals
	wire wrProc31West;
	wire fullProc31West;
	wire [31:0] dataOutProc31West;

	//Processor 32 control and data signals
	wire rdProc32North;
	wire emptyProc32North;
	wire [31:0] dataInProc32North;

	 //Processor 32 control and data signals
	wire wrProc32North;
	wire fullProc32North;
	wire [31:0] dataOutProc32North;

	 //Processor 32 control and data signals
	wire rdProc32South;
	wire emptyProc32South;
	wire [31:0] dataInProc32South;
	
	 //Processor 32 control and data signals
	wire wrProc32South;
	wire fullProc32South;
	wire [31:0] dataOutProc32South;

	 //Processor 32 control and data signals
	wire rdProc32East;
	wire emptyProc32East;
	wire [31:0] dataInProc32East;
	
	 //Processor 32 control and data signals
	wire wrProc32East;
	wire fullProc32East;
	wire [31:0] dataOutProc32East;

	 //Processor 32 control and data signals
	wire rdProc32West;
	wire emptyProc32West;
	wire [31:0] dataInProc32West;

	 //Processor 32 control and data signals
	wire wrProc32West;
	wire fullProc32West;
	wire [31:0] dataOutProc32West;

	//Processor 33 control and data signals
	wire rdProc33North;
	wire emptyProc33North;
	wire [31:0] dataInProc33North;

	 //Processor 33 control and data signals
	wire wrProc33North;
	wire fullProc33North;
	wire [31:0] dataOutProc33North;

	 //Processor 33 control and data signals
	wire rdProc33South;
	wire emptyProc33South;
	wire [31:0] dataInProc33South;
	
	 //Processor 33 control and data signals
	wire wrProc33South;
	wire fullProc33South;
	wire [31:0] dataOutProc33South;

	 //Processor 33 control and data signals
	wire rdProc33East;
	wire emptyProc33East;
	wire [31:0] dataInProc33East;
	
	 //Processor 33 control and data signals
	wire wrProc33East;
	wire fullProc33East;
	wire [31:0] dataOutProc33East;

	 //Processor 33 control and data signals
	wire rdProc33West;
	wire emptyProc33West;
	wire [31:0] dataInProc33West;

	 //Processor 33 control and data signals
	wire wrProc33West;
	wire fullProc33West;
	wire [31:0] dataOutProc33West;

	//Processor 34 control and data signals
	wire rdProc34North;
	wire emptyProc34North;
	wire [31:0] dataInProc34North;

	 //Processor 34 control and data signals
	wire wrProc34North;
	wire fullProc34North;
	wire [31:0] dataOutProc34North;

	 //Processor 34 control and data signals
	wire rdProc34South;
	wire emptyProc34South;
	wire [31:0] dataInProc34South;
	
	 //Processor 34 control and data signals
	wire wrProc34South;
	wire fullProc34South;
	wire [31:0] dataOutProc34South;

	 //Processor 34 control and data signals
	wire rdProc34East;
	wire emptyProc34East;
	wire [31:0] dataInProc34East;
	
	 //Processor 34 control and data signals
	wire wrProc34East;
	wire fullProc34East;
	wire [31:0] dataOutProc34East;

	 //Processor 34 control and data signals
	wire rdProc34West;
	wire emptyProc34West;
	wire [31:0] dataInProc34West;

	 //Processor 34 control and data signals
	wire wrProc34West;
	wire fullProc34West;
	wire [31:0] dataOutProc34West;

	//Processor 35 control and data signals
	wire rdProc35North;
	wire emptyProc35North;
	wire [31:0] dataInProc35North;

	 //Processor 35 control and data signals
	wire wrProc35North;
	wire fullProc35North;
	wire [31:0] dataOutProc35North;

	 //Processor 35 control and data signals
	wire rdProc35South;
	wire emptyProc35South;
	wire [31:0] dataInProc35South;
	
	 //Processor 35 control and data signals
	wire wrProc35South;
	wire fullProc35South;
	wire [31:0] dataOutProc35South;

	 //Processor 35 control and data signals
	wire rdProc35East;
	wire emptyProc35East;
	wire [31:0] dataInProc35East;
	
	 //Processor 35 control and data signals
	wire wrProc35East;
	wire fullProc35East;
	wire [31:0] dataOutProc35East;

	 //Processor 35 control and data signals
	wire rdProc35West;
	wire emptyProc35West;
	wire [31:0] dataInProc35West;

	 //Processor 35 control and data signals
	wire wrProc35West;
	wire fullProc35West;
	wire [31:0] dataOutProc35West;

	//Processor 36 control and data signals
	wire rdProc36North;
	wire emptyProc36North;
	wire [31:0] dataInProc36North;

	 //Processor 36 control and data signals
	wire wrProc36North;
	wire fullProc36North;
	wire [31:0] dataOutProc36North;

	 //Processor 36 control and data signals
	wire rdProc36South;
	wire emptyProc36South;
	wire [31:0] dataInProc36South;
	
	 //Processor 36 control and data signals
	wire wrProc36South;
	wire fullProc36South;
	wire [31:0] dataOutProc36South;

	 //Processor 36 control and data signals
	wire rdProc36East;
	wire emptyProc36East;
	wire [31:0] dataInProc36East;
	
	 //Processor 36 control and data signals
	wire wrProc36East;
	wire fullProc36East;
	wire [31:0] dataOutProc36East;

	 //Processor 36 control and data signals
	wire rdProc36West;
	wire emptyProc36West;
	wire [31:0] dataInProc36West;

	 //Processor 36 control and data signals
	wire wrProc36West;
	wire fullProc36West;
	wire [31:0] dataOutProc36West;

	//Processor 37 control and data signals
	wire rdProc37North;
	wire emptyProc37North;
	wire [31:0] dataInProc37North;

	 //Processor 37 control and data signals
	wire wrProc37North;
	wire fullProc37North;
	wire [31:0] dataOutProc37North;

	 //Processor 37 control and data signals
	wire rdProc37South;
	wire emptyProc37South;
	wire [31:0] dataInProc37South;
	
	 //Processor 37 control and data signals
	wire wrProc37South;
	wire fullProc37South;
	wire [31:0] dataOutProc37South;

	 //Processor 37 control and data signals
	wire rdProc37East;
	wire emptyProc37East;
	wire [31:0] dataInProc37East;
	
	 //Processor 37 control and data signals
	wire wrProc37East;
	wire fullProc37East;
	wire [31:0] dataOutProc37East;

	 //Processor 37 control and data signals
	wire rdProc37West;
	wire emptyProc37West;
	wire [31:0] dataInProc37West;

	 //Processor 37 control and data signals
	wire wrProc37West;
	wire fullProc37West;
	wire [31:0] dataOutProc37West;

	//Processor 38 control and data signals
	wire wrProc38North;
	wire fullProc38North;
	wire [31:0] dataOutProc38North;

	//Processor 38 control and data signals
        wire rdProc38North;
        wire emptyProc38North;
        wire [31:0] dataInProc38North;

	//Processor 38 control and data signals
	wire rdProc38South;
	wire emptyProc38South;
	wire [31:0] dataInProc38South;
		
	 //Processor 38 control and data signals
	wire wrProc38South;
	wire fullProc38South;
	wire [31:0] dataOutProc38South;

	 //Processor 38 control and data signals
	wire wrProc38West;
	wire fullProc38West;
	wire [31:0] dataOutProc38West;
	
	 //Processor 38 control and data signals
	wire rdProc38West;
	wire emptyProc38West;
	wire [31:0] dataInProc38West;

	//Processor 39 control and data signals
	wire wrProc39North;
	wire fullProc39North;
	wire [31:0] dataOutProc39North;

	 //Processor 39 control and data signals
	wire rdProc39North;
	wire emptyProc39North;
	wire [31:0] dataInProc39North;
	
	 //Processor 39 control and data signals
	wire rdProc39South;
	wire emptyProc39South;
	wire [31:0] dataInProc39South;
	
	 //Processor 39 control and data signals
	wire wrProc39South;
	wire fullProc39South;
	wire [31:0] dataOutProc39South;
	
	 //Processor 39 control and data signals
	wire rdProc39East;
	wire emptyProc39East;
	wire [31:0] dataInProc39East;

	 //Processor 39 control and data signals
	wire wrProc39East;
	wire fullProc39East;
	wire [31:0] dataOutProc39East;

	//Processor 40 control and data signals
	wire rdProc40North;
	wire emptyProc40North;
	wire [31:0] dataInProc40North;

	 //Processor 40 control and data signals
	wire wrProc40North;
	wire fullProc40North;
	wire [31:0] dataOutProc40North;

	 //Processor 40 control and data signals
	wire rdProc40South;
	wire emptyProc40South;
	wire [31:0] dataInProc40South;
	
	 //Processor 40 control and data signals
	wire wrProc40South;
	wire fullProc40South;
	wire [31:0] dataOutProc40South;

	 //Processor 40 control and data signals
	wire rdProc40East;
	wire emptyProc40East;
	wire [31:0] dataInProc40East;
	
	 //Processor 40 control and data signals
	wire wrProc40East;
	wire fullProc40East;
	wire [31:0] dataOutProc40East;

	 //Processor 40 control and data signals
	wire rdProc40West;
	wire emptyProc40West;
	wire [31:0] dataInProc40West;

	 //Processor 40 control and data signals
	wire wrProc40West;
	wire fullProc40West;
	wire [31:0] dataOutProc40West;

	//Processor 41 control and data signals
	wire rdProc41North;
	wire emptyProc41North;
	wire [31:0] dataInProc41North;

	 //Processor 41 control and data signals
	wire wrProc41North;
	wire fullProc41North;
	wire [31:0] dataOutProc41North;

	 //Processor 41 control and data signals
	wire rdProc41South;
	wire emptyProc41South;
	wire [31:0] dataInProc41South;
	
	 //Processor 41 control and data signals
	wire wrProc41South;
	wire fullProc41South;
	wire [31:0] dataOutProc41South;

	 //Processor 41 control and data signals
	wire rdProc41East;
	wire emptyProc41East;
	wire [31:0] dataInProc41East;
	
	 //Processor 41 control and data signals
	wire wrProc41East;
	wire fullProc41East;
	wire [31:0] dataOutProc41East;

	 //Processor 41 control and data signals
	wire rdProc41West;
	wire emptyProc41West;
	wire [31:0] dataInProc41West;

	 //Processor 41 control and data signals
	wire wrProc41West;
	wire fullProc41West;
	wire [31:0] dataOutProc41West;

	//Processor 42 control and data signals
	wire rdProc42North;
	wire emptyProc42North;
	wire [31:0] dataInProc42North;

	 //Processor 42 control and data signals
	wire wrProc42North;
	wire fullProc42North;
	wire [31:0] dataOutProc42North;

	 //Processor 42 control and data signals
	wire rdProc42South;
	wire emptyProc42South;
	wire [31:0] dataInProc42South;
	
	 //Processor 42 control and data signals
	wire wrProc42South;
	wire fullProc42South;
	wire [31:0] dataOutProc42South;

	 //Processor 42 control and data signals
	wire rdProc42East;
	wire emptyProc42East;
	wire [31:0] dataInProc42East;
	
	 //Processor 42 control and data signals
	wire wrProc42East;
	wire fullProc42East;
	wire [31:0] dataOutProc42East;

	 //Processor 42 control and data signals
	wire rdProc42West;
	wire emptyProc42West;
	wire [31:0] dataInProc42West;

	 //Processor 42 control and data signals
	wire wrProc42West;
	wire fullProc42West;
	wire [31:0] dataOutProc42West;

	//Processor 43 control and data signals
	wire rdProc43North;
	wire emptyProc43North;
	wire [31:0] dataInProc43North;

	 //Processor 43 control and data signals
	wire wrProc43North;
	wire fullProc43North;
	wire [31:0] dataOutProc43North;

	 //Processor 43 control and data signals
	wire rdProc43South;
	wire emptyProc43South;
	wire [31:0] dataInProc43South;
	
	 //Processor 43 control and data signals
	wire wrProc43South;
	wire fullProc43South;
	wire [31:0] dataOutProc43South;

	 //Processor 43 control and data signals
	wire rdProc43East;
	wire emptyProc43East;
	wire [31:0] dataInProc43East;
	
	 //Processor 43 control and data signals
	wire wrProc43East;
	wire fullProc43East;
	wire [31:0] dataOutProc43East;

	 //Processor 43 control and data signals
	wire rdProc43West;
	wire emptyProc43West;
	wire [31:0] dataInProc43West;

	 //Processor 43 control and data signals
	wire wrProc43West;
	wire fullProc43West;
	wire [31:0] dataOutProc43West;

	//Processor 44 control and data signals
	wire rdProc44North;
	wire emptyProc44North;
	wire [31:0] dataInProc44North;

	 //Processor 44 control and data signals
	wire wrProc44North;
	wire fullProc44North;
	wire [31:0] dataOutProc44North;

	 //Processor 44 control and data signals
	wire rdProc44South;
	wire emptyProc44South;
	wire [31:0] dataInProc44South;
	
	 //Processor 44 control and data signals
	wire wrProc44South;
	wire fullProc44South;
	wire [31:0] dataOutProc44South;

	 //Processor 44 control and data signals
	wire rdProc44East;
	wire emptyProc44East;
	wire [31:0] dataInProc44East;
	
	 //Processor 44 control and data signals
	wire wrProc44East;
	wire fullProc44East;
	wire [31:0] dataOutProc44East;

	 //Processor 44 control and data signals
	wire rdProc44West;
	wire emptyProc44West;
	wire [31:0] dataInProc44West;

	 //Processor 44 control and data signals
	wire wrProc44West;
	wire fullProc44West;
	wire [31:0] dataOutProc44West;

	//Processor 45 control and data signals
	wire rdProc45North;
	wire emptyProc45North;
	wire [31:0] dataInProc45North;

	 //Processor 45 control and data signals
	wire wrProc45North;
	wire fullProc45North;
	wire [31:0] dataOutProc45North;

	 //Processor 45 control and data signals
	wire rdProc45South;
	wire emptyProc45South;
	wire [31:0] dataInProc45South;
	
	 //Processor 45 control and data signals
	wire wrProc45South;
	wire fullProc45South;
	wire [31:0] dataOutProc45South;

	 //Processor 45 control and data signals
	wire rdProc45East;
	wire emptyProc45East;
	wire [31:0] dataInProc45East;
	
	 //Processor 45 control and data signals
	wire wrProc45East;
	wire fullProc45East;
	wire [31:0] dataOutProc45East;

	 //Processor 45 control and data signals
	wire rdProc45West;
	wire emptyProc45West;
	wire [31:0] dataInProc45West;

	 //Processor 45 control and data signals
	wire wrProc45West;
	wire fullProc45West;
	wire [31:0] dataOutProc45West;

	//Processor 46 control and data signals
	wire rdProc46North;
	wire emptyProc46North;
	wire [31:0] dataInProc46North;

	 //Processor 46 control and data signals
	wire wrProc46North;
	wire fullProc46North;
	wire [31:0] dataOutProc46North;

	 //Processor 46 control and data signals
	wire rdProc46South;
	wire emptyProc46South;
	wire [31:0] dataInProc46South;
	
	 //Processor 46 control and data signals
	wire wrProc46South;
	wire fullProc46South;
	wire [31:0] dataOutProc46South;

	 //Processor 46 control and data signals
	wire rdProc46East;
	wire emptyProc46East;
	wire [31:0] dataInProc46East;
	
	 //Processor 46 control and data signals
	wire wrProc46East;
	wire fullProc46East;
	wire [31:0] dataOutProc46East;

	 //Processor 46 control and data signals
	wire rdProc46West;
	wire emptyProc46West;
	wire [31:0] dataInProc46West;

	 //Processor 46 control and data signals
	wire wrProc46West;
	wire fullProc46West;
	wire [31:0] dataOutProc46West;

	//Processor 47 control and data signals
	wire rdProc47North;
	wire emptyProc47North;
	wire [31:0] dataInProc47North;

	 //Processor 47 control and data signals
	wire wrProc47North;
	wire fullProc47North;
	wire [31:0] dataOutProc47North;

	 //Processor 47 control and data signals
	wire rdProc47South;
	wire emptyProc47South;
	wire [31:0] dataInProc47South;
	
	 //Processor 47 control and data signals
	wire wrProc47South;
	wire fullProc47South;
	wire [31:0] dataOutProc47South;

	 //Processor 47 control and data signals
	wire rdProc47East;
	wire emptyProc47East;
	wire [31:0] dataInProc47East;
	
	 //Processor 47 control and data signals
	wire wrProc47East;
	wire fullProc47East;
	wire [31:0] dataOutProc47East;

	 //Processor 47 control and data signals
	wire rdProc47West;
	wire emptyProc47West;
	wire [31:0] dataInProc47West;

	 //Processor 47 control and data signals
	wire wrProc47West;
	wire fullProc47West;
	wire [31:0] dataOutProc47West;

	//Processor 48 control and data signals
	wire rdProc48North;
	wire emptyProc48North;
	wire [31:0] dataInProc48North;

	 //Processor 48 control and data signals
	wire wrProc48North;
	wire fullProc48North;
	wire [31:0] dataOutProc48North;

	 //Processor 48 control and data signals
	wire rdProc48South;
	wire emptyProc48South;
	wire [31:0] dataInProc48South;
	
	 //Processor 48 control and data signals
	wire wrProc48South;
	wire fullProc48South;
	wire [31:0] dataOutProc48South;

	 //Processor 48 control and data signals
	wire rdProc48East;
	wire emptyProc48East;
	wire [31:0] dataInProc48East;
	
	 //Processor 48 control and data signals
	wire wrProc48East;
	wire fullProc48East;
	wire [31:0] dataOutProc48East;

	 //Processor 48 control and data signals
	wire rdProc48West;
	wire emptyProc48West;
	wire [31:0] dataInProc48West;

	 //Processor 48 control and data signals
	wire wrProc48West;
	wire fullProc48West;
	wire [31:0] dataOutProc48West;

	//Processor 49 control and data signals
	wire rdProc49North;
	wire emptyProc49North;
	wire [31:0] dataInProc49North;

	 //Processor 49 control and data signals
	wire wrProc49North;
	wire fullProc49North;
	wire [31:0] dataOutProc49North;

	 //Processor 49 control and data signals
	wire rdProc49South;
	wire emptyProc49South;
	wire [31:0] dataInProc49South;
	
	 //Processor 49 control and data signals
	wire wrProc49South;
	wire fullProc49South;
	wire [31:0] dataOutProc49South;

	 //Processor 49 control and data signals
	wire rdProc49East;
	wire emptyProc49East;
	wire [31:0] dataInProc49East;
	
	 //Processor 49 control and data signals
	wire wrProc49East;
	wire fullProc49East;
	wire [31:0] dataOutProc49East;

	 //Processor 49 control and data signals
	wire rdProc49West;
	wire emptyProc49West;
	wire [31:0] dataInProc49West;

	 //Processor 49 control and data signals
	wire wrProc49West;
	wire fullProc49West;
	wire [31:0] dataOutProc49West;

	//Processor 50 control and data signals
	wire rdProc50North;
	wire emptyProc50North;
	wire [31:0] dataInProc50North;

	 //Processor 50 control and data signals
	wire wrProc50North;
	wire fullProc50North;
	wire [31:0] dataOutProc50North;

	 //Processor 50 control and data signals
	wire rdProc50South;
	wire emptyProc50South;
	wire [31:0] dataInProc50South;
	
	 //Processor 50 control and data signals
	wire wrProc50South;
	wire fullProc50South;
	wire [31:0] dataOutProc50South;

	 //Processor 50 control and data signals
	wire rdProc50East;
	wire emptyProc50East;
	wire [31:0] dataInProc50East;
	
	 //Processor 50 control and data signals
	wire wrProc50East;
	wire fullProc50East;
	wire [31:0] dataOutProc50East;

	 //Processor 50 control and data signals
	wire rdProc50West;
	wire emptyProc50West;
	wire [31:0] dataInProc50West;

	 //Processor 50 control and data signals
	wire wrProc50West;
	wire fullProc50West;
	wire [31:0] dataOutProc50West;

	//Processor 51 control and data signals
	wire wrProc51North;
	wire fullProc51North;
	wire [31:0] dataOutProc51North;

	//Processor 51 control and data signals
        wire rdProc51North;
        wire emptyProc51North;
        wire [31:0] dataInProc51North;

	//Processor 51 control and data signals
	wire rdProc51South;
	wire emptyProc51South;
	wire [31:0] dataInProc51South;
		
	 //Processor 51 control and data signals
	wire wrProc51South;
	wire fullProc51South;
	wire [31:0] dataOutProc51South;

	 //Processor 51 control and data signals
	wire wrProc51West;
	wire fullProc51West;
	wire [31:0] dataOutProc51West;
	
	 //Processor 51 control and data signals
	wire rdProc51West;
	wire emptyProc51West;
	wire [31:0] dataInProc51West;

	//Processor 52 control and data signals
	wire wrProc52North;
	wire fullProc52North;
	wire [31:0] dataOutProc52North;

	 //Processor 52 control and data signals
	wire rdProc52North;
	wire emptyProc52North;
	wire [31:0] dataInProc52North;
	
	 //Processor 52 control and data signals
	wire rdProc52South;
	wire emptyProc52South;
	wire [31:0] dataInProc52South;
	
	 //Processor 52 control and data signals
	wire wrProc52South;
	wire fullProc52South;
	wire [31:0] dataOutProc52South;
	
	 //Processor 52 control and data signals
	wire rdProc52East;
	wire emptyProc52East;
	wire [31:0] dataInProc52East;

	 //Processor 52 control and data signals
	wire wrProc52East;
	wire fullProc52East;
	wire [31:0] dataOutProc52East;

	//Processor 53 control and data signals
	wire rdProc53North;
	wire emptyProc53North;
	wire [31:0] dataInProc53North;

	 //Processor 53 control and data signals
	wire wrProc53North;
	wire fullProc53North;
	wire [31:0] dataOutProc53North;

	 //Processor 53 control and data signals
	wire rdProc53South;
	wire emptyProc53South;
	wire [31:0] dataInProc53South;
	
	 //Processor 53 control and data signals
	wire wrProc53South;
	wire fullProc53South;
	wire [31:0] dataOutProc53South;

	 //Processor 53 control and data signals
	wire rdProc53East;
	wire emptyProc53East;
	wire [31:0] dataInProc53East;
	
	 //Processor 53 control and data signals
	wire wrProc53East;
	wire fullProc53East;
	wire [31:0] dataOutProc53East;

	 //Processor 53 control and data signals
	wire rdProc53West;
	wire emptyProc53West;
	wire [31:0] dataInProc53West;

	 //Processor 53 control and data signals
	wire wrProc53West;
	wire fullProc53West;
	wire [31:0] dataOutProc53West;

	//Processor 54 control and data signals
	wire rdProc54North;
	wire emptyProc54North;
	wire [31:0] dataInProc54North;

	 //Processor 54 control and data signals
	wire wrProc54North;
	wire fullProc54North;
	wire [31:0] dataOutProc54North;

	 //Processor 54 control and data signals
	wire rdProc54South;
	wire emptyProc54South;
	wire [31:0] dataInProc54South;
	
	 //Processor 54 control and data signals
	wire wrProc54South;
	wire fullProc54South;
	wire [31:0] dataOutProc54South;

	 //Processor 54 control and data signals
	wire rdProc54East;
	wire emptyProc54East;
	wire [31:0] dataInProc54East;
	
	 //Processor 54 control and data signals
	wire wrProc54East;
	wire fullProc54East;
	wire [31:0] dataOutProc54East;

	 //Processor 54 control and data signals
	wire rdProc54West;
	wire emptyProc54West;
	wire [31:0] dataInProc54West;

	 //Processor 54 control and data signals
	wire wrProc54West;
	wire fullProc54West;
	wire [31:0] dataOutProc54West;

	//Processor 55 control and data signals
	wire rdProc55North;
	wire emptyProc55North;
	wire [31:0] dataInProc55North;

	 //Processor 55 control and data signals
	wire wrProc55North;
	wire fullProc55North;
	wire [31:0] dataOutProc55North;

	 //Processor 55 control and data signals
	wire rdProc55South;
	wire emptyProc55South;
	wire [31:0] dataInProc55South;
	
	 //Processor 55 control and data signals
	wire wrProc55South;
	wire fullProc55South;
	wire [31:0] dataOutProc55South;

	 //Processor 55 control and data signals
	wire rdProc55East;
	wire emptyProc55East;
	wire [31:0] dataInProc55East;
	
	 //Processor 55 control and data signals
	wire wrProc55East;
	wire fullProc55East;
	wire [31:0] dataOutProc55East;

	 //Processor 55 control and data signals
	wire rdProc55West;
	wire emptyProc55West;
	wire [31:0] dataInProc55West;

	 //Processor 55 control and data signals
	wire wrProc55West;
	wire fullProc55West;
	wire [31:0] dataOutProc55West;

	//Processor 56 control and data signals
	wire rdProc56North;
	wire emptyProc56North;
	wire [31:0] dataInProc56North;

	 //Processor 56 control and data signals
	wire wrProc56North;
	wire fullProc56North;
	wire [31:0] dataOutProc56North;

	 //Processor 56 control and data signals
	wire rdProc56South;
	wire emptyProc56South;
	wire [31:0] dataInProc56South;
	
	 //Processor 56 control and data signals
	wire wrProc56South;
	wire fullProc56South;
	wire [31:0] dataOutProc56South;

	 //Processor 56 control and data signals
	wire rdProc56East;
	wire emptyProc56East;
	wire [31:0] dataInProc56East;
	
	 //Processor 56 control and data signals
	wire wrProc56East;
	wire fullProc56East;
	wire [31:0] dataOutProc56East;

	 //Processor 56 control and data signals
	wire rdProc56West;
	wire emptyProc56West;
	wire [31:0] dataInProc56West;

	 //Processor 56 control and data signals
	wire wrProc56West;
	wire fullProc56West;
	wire [31:0] dataOutProc56West;

	//Processor 57 control and data signals
	wire rdProc57North;
	wire emptyProc57North;
	wire [31:0] dataInProc57North;

	 //Processor 57 control and data signals
	wire wrProc57North;
	wire fullProc57North;
	wire [31:0] dataOutProc57North;

	 //Processor 57 control and data signals
	wire rdProc57South;
	wire emptyProc57South;
	wire [31:0] dataInProc57South;
	
	 //Processor 57 control and data signals
	wire wrProc57South;
	wire fullProc57South;
	wire [31:0] dataOutProc57South;

	 //Processor 57 control and data signals
	wire rdProc57East;
	wire emptyProc57East;
	wire [31:0] dataInProc57East;
	
	 //Processor 57 control and data signals
	wire wrProc57East;
	wire fullProc57East;
	wire [31:0] dataOutProc57East;

	 //Processor 57 control and data signals
	wire rdProc57West;
	wire emptyProc57West;
	wire [31:0] dataInProc57West;

	 //Processor 57 control and data signals
	wire wrProc57West;
	wire fullProc57West;
	wire [31:0] dataOutProc57West;

	//Processor 58 control and data signals
	wire rdProc58North;
	wire emptyProc58North;
	wire [31:0] dataInProc58North;

	 //Processor 58 control and data signals
	wire wrProc58North;
	wire fullProc58North;
	wire [31:0] dataOutProc58North;

	 //Processor 58 control and data signals
	wire rdProc58South;
	wire emptyProc58South;
	wire [31:0] dataInProc58South;
	
	 //Processor 58 control and data signals
	wire wrProc58South;
	wire fullProc58South;
	wire [31:0] dataOutProc58South;

	 //Processor 58 control and data signals
	wire rdProc58East;
	wire emptyProc58East;
	wire [31:0] dataInProc58East;
	
	 //Processor 58 control and data signals
	wire wrProc58East;
	wire fullProc58East;
	wire [31:0] dataOutProc58East;

	 //Processor 58 control and data signals
	wire rdProc58West;
	wire emptyProc58West;
	wire [31:0] dataInProc58West;

	 //Processor 58 control and data signals
	wire wrProc58West;
	wire fullProc58West;
	wire [31:0] dataOutProc58West;

	//Processor 59 control and data signals
	wire rdProc59North;
	wire emptyProc59North;
	wire [31:0] dataInProc59North;

	 //Processor 59 control and data signals
	wire wrProc59North;
	wire fullProc59North;
	wire [31:0] dataOutProc59North;

	 //Processor 59 control and data signals
	wire rdProc59South;
	wire emptyProc59South;
	wire [31:0] dataInProc59South;
	
	 //Processor 59 control and data signals
	wire wrProc59South;
	wire fullProc59South;
	wire [31:0] dataOutProc59South;

	 //Processor 59 control and data signals
	wire rdProc59East;
	wire emptyProc59East;
	wire [31:0] dataInProc59East;
	
	 //Processor 59 control and data signals
	wire wrProc59East;
	wire fullProc59East;
	wire [31:0] dataOutProc59East;

	 //Processor 59 control and data signals
	wire rdProc59West;
	wire emptyProc59West;
	wire [31:0] dataInProc59West;

	 //Processor 59 control and data signals
	wire wrProc59West;
	wire fullProc59West;
	wire [31:0] dataOutProc59West;

	//Processor 60 control and data signals
	wire rdProc60North;
	wire emptyProc60North;
	wire [31:0] dataInProc60North;

	 //Processor 60 control and data signals
	wire wrProc60North;
	wire fullProc60North;
	wire [31:0] dataOutProc60North;

	 //Processor 60 control and data signals
	wire rdProc60South;
	wire emptyProc60South;
	wire [31:0] dataInProc60South;
	
	 //Processor 60 control and data signals
	wire wrProc60South;
	wire fullProc60South;
	wire [31:0] dataOutProc60South;

	 //Processor 60 control and data signals
	wire rdProc60East;
	wire emptyProc60East;
	wire [31:0] dataInProc60East;
	
	 //Processor 60 control and data signals
	wire wrProc60East;
	wire fullProc60East;
	wire [31:0] dataOutProc60East;

	 //Processor 60 control and data signals
	wire rdProc60West;
	wire emptyProc60West;
	wire [31:0] dataInProc60West;

	 //Processor 60 control and data signals
	wire wrProc60West;
	wire fullProc60West;
	wire [31:0] dataOutProc60West;

	//Processor 61 control and data signals
	wire rdProc61North;
	wire emptyProc61North;
	wire [31:0] dataInProc61North;

	 //Processor 61 control and data signals
	wire wrProc61North;
	wire fullProc61North;
	wire [31:0] dataOutProc61North;

	 //Processor 61 control and data signals
	wire rdProc61South;
	wire emptyProc61South;
	wire [31:0] dataInProc61South;
	
	 //Processor 61 control and data signals
	wire wrProc61South;
	wire fullProc61South;
	wire [31:0] dataOutProc61South;

	 //Processor 61 control and data signals
	wire rdProc61East;
	wire emptyProc61East;
	wire [31:0] dataInProc61East;
	
	 //Processor 61 control and data signals
	wire wrProc61East;
	wire fullProc61East;
	wire [31:0] dataOutProc61East;

	 //Processor 61 control and data signals
	wire rdProc61West;
	wire emptyProc61West;
	wire [31:0] dataInProc61West;

	 //Processor 61 control and data signals
	wire wrProc61West;
	wire fullProc61West;
	wire [31:0] dataOutProc61West;

	//Processor 62 control and data signals
	wire rdProc62North;
	wire emptyProc62North;
	wire [31:0] dataInProc62North;

	 //Processor 62 control and data signals
	wire wrProc62North;
	wire fullProc62North;
	wire [31:0] dataOutProc62North;

	 //Processor 62 control and data signals
	wire rdProc62South;
	wire emptyProc62South;
	wire [31:0] dataInProc62South;
	
	 //Processor 62 control and data signals
	wire wrProc62South;
	wire fullProc62South;
	wire [31:0] dataOutProc62South;

	 //Processor 62 control and data signals
	wire rdProc62East;
	wire emptyProc62East;
	wire [31:0] dataInProc62East;
	
	 //Processor 62 control and data signals
	wire wrProc62East;
	wire fullProc62East;
	wire [31:0] dataOutProc62East;

	 //Processor 62 control and data signals
	wire rdProc62West;
	wire emptyProc62West;
	wire [31:0] dataInProc62West;

	 //Processor 62 control and data signals
	wire wrProc62West;
	wire fullProc62West;
	wire [31:0] dataOutProc62West;

	//Processor 63 control and data signals
	wire rdProc63North;
	wire emptyProc63North;
	wire [31:0] dataInProc63North;

	 //Processor 63 control and data signals
	wire wrProc63North;
	wire fullProc63North;
	wire [31:0] dataOutProc63North;

	 //Processor 63 control and data signals
	wire rdProc63South;
	wire emptyProc63South;
	wire [31:0] dataInProc63South;
	
	 //Processor 63 control and data signals
	wire wrProc63South;
	wire fullProc63South;
	wire [31:0] dataOutProc63South;

	 //Processor 63 control and data signals
	wire rdProc63East;
	wire emptyProc63East;
	wire [31:0] dataInProc63East;
	
	 //Processor 63 control and data signals
	wire wrProc63East;
	wire fullProc63East;
	wire [31:0] dataOutProc63East;

	 //Processor 63 control and data signals
	wire rdProc63West;
	wire emptyProc63West;
	wire [31:0] dataInProc63West;

	 //Processor 63 control and data signals
	wire wrProc63West;
	wire fullProc63West;
	wire [31:0] dataOutProc63West;

	//Processor 64 control and data signals
	wire wrProc64North;
	wire fullProc64North;
	wire [31:0] dataOutProc64North;

	//Processor 64 control and data signals
        wire rdProc64North;
        wire emptyProc64North;
        wire [31:0] dataInProc64North;

	//Processor 64 control and data signals
	wire rdProc64South;
	wire emptyProc64South;
	wire [31:0] dataInProc64South;
		
	 //Processor 64 control and data signals
	wire wrProc64South;
	wire fullProc64South;
	wire [31:0] dataOutProc64South;

	 //Processor 64 control and data signals
	wire wrProc64West;
	wire fullProc64West;
	wire [31:0] dataOutProc64West;
	
	 //Processor 64 control and data signals
	wire rdProc64West;
	wire emptyProc64West;
	wire [31:0] dataInProc64West;

	//Processor 65 control and data signals
	wire wrProc65North;
	wire fullProc65North;
	wire [31:0] dataOutProc65North;

	 //Processor 65 control and data signals
	wire rdProc65North;
	wire emptyProc65North;
	wire [31:0] dataInProc65North;
	
	 //Processor 65 control and data signals
	wire rdProc65South;
	wire emptyProc65South;
	wire [31:0] dataInProc65South;
	
	 //Processor 65 control and data signals
	wire wrProc65South;
	wire fullProc65South;
	wire [31:0] dataOutProc65South;
	
	 //Processor 65 control and data signals
	wire rdProc65East;
	wire emptyProc65East;
	wire [31:0] dataInProc65East;

	 //Processor 65 control and data signals
	wire wrProc65East;
	wire fullProc65East;
	wire [31:0] dataOutProc65East;

	//Processor 66 control and data signals
	wire rdProc66North;
	wire emptyProc66North;
	wire [31:0] dataInProc66North;

	 //Processor 66 control and data signals
	wire wrProc66North;
	wire fullProc66North;
	wire [31:0] dataOutProc66North;

	 //Processor 66 control and data signals
	wire rdProc66South;
	wire emptyProc66South;
	wire [31:0] dataInProc66South;
	
	 //Processor 66 control and data signals
	wire wrProc66South;
	wire fullProc66South;
	wire [31:0] dataOutProc66South;

	 //Processor 66 control and data signals
	wire rdProc66East;
	wire emptyProc66East;
	wire [31:0] dataInProc66East;
	
	 //Processor 66 control and data signals
	wire wrProc66East;
	wire fullProc66East;
	wire [31:0] dataOutProc66East;

	 //Processor 66 control and data signals
	wire rdProc66West;
	wire emptyProc66West;
	wire [31:0] dataInProc66West;

	 //Processor 66 control and data signals
	wire wrProc66West;
	wire fullProc66West;
	wire [31:0] dataOutProc66West;

	//Processor 67 control and data signals
	wire rdProc67North;
	wire emptyProc67North;
	wire [31:0] dataInProc67North;

	 //Processor 67 control and data signals
	wire wrProc67North;
	wire fullProc67North;
	wire [31:0] dataOutProc67North;

	 //Processor 67 control and data signals
	wire rdProc67South;
	wire emptyProc67South;
	wire [31:0] dataInProc67South;
	
	 //Processor 67 control and data signals
	wire wrProc67South;
	wire fullProc67South;
	wire [31:0] dataOutProc67South;

	 //Processor 67 control and data signals
	wire rdProc67East;
	wire emptyProc67East;
	wire [31:0] dataInProc67East;
	
	 //Processor 67 control and data signals
	wire wrProc67East;
	wire fullProc67East;
	wire [31:0] dataOutProc67East;

	 //Processor 67 control and data signals
	wire rdProc67West;
	wire emptyProc67West;
	wire [31:0] dataInProc67West;

	 //Processor 67 control and data signals
	wire wrProc67West;
	wire fullProc67West;
	wire [31:0] dataOutProc67West;

	//Processor 68 control and data signals
	wire rdProc68North;
	wire emptyProc68North;
	wire [31:0] dataInProc68North;

	 //Processor 68 control and data signals
	wire wrProc68North;
	wire fullProc68North;
	wire [31:0] dataOutProc68North;

	 //Processor 68 control and data signals
	wire rdProc68South;
	wire emptyProc68South;
	wire [31:0] dataInProc68South;
	
	 //Processor 68 control and data signals
	wire wrProc68South;
	wire fullProc68South;
	wire [31:0] dataOutProc68South;

	 //Processor 68 control and data signals
	wire rdProc68East;
	wire emptyProc68East;
	wire [31:0] dataInProc68East;
	
	 //Processor 68 control and data signals
	wire wrProc68East;
	wire fullProc68East;
	wire [31:0] dataOutProc68East;

	 //Processor 68 control and data signals
	wire rdProc68West;
	wire emptyProc68West;
	wire [31:0] dataInProc68West;

	 //Processor 68 control and data signals
	wire wrProc68West;
	wire fullProc68West;
	wire [31:0] dataOutProc68West;

	//Processor 69 control and data signals
	wire rdProc69North;
	wire emptyProc69North;
	wire [31:0] dataInProc69North;

	 //Processor 69 control and data signals
	wire wrProc69North;
	wire fullProc69North;
	wire [31:0] dataOutProc69North;

	 //Processor 69 control and data signals
	wire rdProc69South;
	wire emptyProc69South;
	wire [31:0] dataInProc69South;
	
	 //Processor 69 control and data signals
	wire wrProc69South;
	wire fullProc69South;
	wire [31:0] dataOutProc69South;

	 //Processor 69 control and data signals
	wire rdProc69East;
	wire emptyProc69East;
	wire [31:0] dataInProc69East;
	
	 //Processor 69 control and data signals
	wire wrProc69East;
	wire fullProc69East;
	wire [31:0] dataOutProc69East;

	 //Processor 69 control and data signals
	wire rdProc69West;
	wire emptyProc69West;
	wire [31:0] dataInProc69West;

	 //Processor 69 control and data signals
	wire wrProc69West;
	wire fullProc69West;
	wire [31:0] dataOutProc69West;

	//Processor 70 control and data signals
	wire rdProc70North;
	wire emptyProc70North;
	wire [31:0] dataInProc70North;

	 //Processor 70 control and data signals
	wire wrProc70North;
	wire fullProc70North;
	wire [31:0] dataOutProc70North;

	 //Processor 70 control and data signals
	wire rdProc70South;
	wire emptyProc70South;
	wire [31:0] dataInProc70South;
	
	 //Processor 70 control and data signals
	wire wrProc70South;
	wire fullProc70South;
	wire [31:0] dataOutProc70South;

	 //Processor 70 control and data signals
	wire rdProc70East;
	wire emptyProc70East;
	wire [31:0] dataInProc70East;
	
	 //Processor 70 control and data signals
	wire wrProc70East;
	wire fullProc70East;
	wire [31:0] dataOutProc70East;

	 //Processor 70 control and data signals
	wire rdProc70West;
	wire emptyProc70West;
	wire [31:0] dataInProc70West;

	 //Processor 70 control and data signals
	wire wrProc70West;
	wire fullProc70West;
	wire [31:0] dataOutProc70West;

	//Processor 71 control and data signals
	wire rdProc71North;
	wire emptyProc71North;
	wire [31:0] dataInProc71North;

	 //Processor 71 control and data signals
	wire wrProc71North;
	wire fullProc71North;
	wire [31:0] dataOutProc71North;

	 //Processor 71 control and data signals
	wire rdProc71South;
	wire emptyProc71South;
	wire [31:0] dataInProc71South;
	
	 //Processor 71 control and data signals
	wire wrProc71South;
	wire fullProc71South;
	wire [31:0] dataOutProc71South;

	 //Processor 71 control and data signals
	wire rdProc71East;
	wire emptyProc71East;
	wire [31:0] dataInProc71East;
	
	 //Processor 71 control and data signals
	wire wrProc71East;
	wire fullProc71East;
	wire [31:0] dataOutProc71East;

	 //Processor 71 control and data signals
	wire rdProc71West;
	wire emptyProc71West;
	wire [31:0] dataInProc71West;

	 //Processor 71 control and data signals
	wire wrProc71West;
	wire fullProc71West;
	wire [31:0] dataOutProc71West;

	//Processor 72 control and data signals
	wire rdProc72North;
	wire emptyProc72North;
	wire [31:0] dataInProc72North;

	 //Processor 72 control and data signals
	wire wrProc72North;
	wire fullProc72North;
	wire [31:0] dataOutProc72North;

	 //Processor 72 control and data signals
	wire rdProc72South;
	wire emptyProc72South;
	wire [31:0] dataInProc72South;
	
	 //Processor 72 control and data signals
	wire wrProc72South;
	wire fullProc72South;
	wire [31:0] dataOutProc72South;

	 //Processor 72 control and data signals
	wire rdProc72East;
	wire emptyProc72East;
	wire [31:0] dataInProc72East;
	
	 //Processor 72 control and data signals
	wire wrProc72East;
	wire fullProc72East;
	wire [31:0] dataOutProc72East;

	 //Processor 72 control and data signals
	wire rdProc72West;
	wire emptyProc72West;
	wire [31:0] dataInProc72West;

	 //Processor 72 control and data signals
	wire wrProc72West;
	wire fullProc72West;
	wire [31:0] dataOutProc72West;

	//Processor 73 control and data signals
	wire rdProc73North;
	wire emptyProc73North;
	wire [31:0] dataInProc73North;

	 //Processor 73 control and data signals
	wire wrProc73North;
	wire fullProc73North;
	wire [31:0] dataOutProc73North;

	 //Processor 73 control and data signals
	wire rdProc73South;
	wire emptyProc73South;
	wire [31:0] dataInProc73South;
	
	 //Processor 73 control and data signals
	wire wrProc73South;
	wire fullProc73South;
	wire [31:0] dataOutProc73South;

	 //Processor 73 control and data signals
	wire rdProc73East;
	wire emptyProc73East;
	wire [31:0] dataInProc73East;
	
	 //Processor 73 control and data signals
	wire wrProc73East;
	wire fullProc73East;
	wire [31:0] dataOutProc73East;

	 //Processor 73 control and data signals
	wire rdProc73West;
	wire emptyProc73West;
	wire [31:0] dataInProc73West;

	 //Processor 73 control and data signals
	wire wrProc73West;
	wire fullProc73West;
	wire [31:0] dataOutProc73West;

	//Processor 74 control and data signals
	wire rdProc74North;
	wire emptyProc74North;
	wire [31:0] dataInProc74North;

	 //Processor 74 control and data signals
	wire wrProc74North;
	wire fullProc74North;
	wire [31:0] dataOutProc74North;

	 //Processor 74 control and data signals
	wire rdProc74South;
	wire emptyProc74South;
	wire [31:0] dataInProc74South;
	
	 //Processor 74 control and data signals
	wire wrProc74South;
	wire fullProc74South;
	wire [31:0] dataOutProc74South;

	 //Processor 74 control and data signals
	wire rdProc74East;
	wire emptyProc74East;
	wire [31:0] dataInProc74East;
	
	 //Processor 74 control and data signals
	wire wrProc74East;
	wire fullProc74East;
	wire [31:0] dataOutProc74East;

	 //Processor 74 control and data signals
	wire rdProc74West;
	wire emptyProc74West;
	wire [31:0] dataInProc74West;

	 //Processor 74 control and data signals
	wire wrProc74West;
	wire fullProc74West;
	wire [31:0] dataOutProc74West;

	//Processor 75 control and data signals
	wire rdProc75North;
	wire emptyProc75North;
	wire [31:0] dataInProc75North;

	 //Processor 75 control and data signals
	wire wrProc75North;
	wire fullProc75North;
	wire [31:0] dataOutProc75North;

	 //Processor 75 control and data signals
	wire rdProc75South;
	wire emptyProc75South;
	wire [31:0] dataInProc75South;
	
	 //Processor 75 control and data signals
	wire wrProc75South;
	wire fullProc75South;
	wire [31:0] dataOutProc75South;

	 //Processor 75 control and data signals
	wire rdProc75East;
	wire emptyProc75East;
	wire [31:0] dataInProc75East;
	
	 //Processor 75 control and data signals
	wire wrProc75East;
	wire fullProc75East;
	wire [31:0] dataOutProc75East;

	 //Processor 75 control and data signals
	wire rdProc75West;
	wire emptyProc75West;
	wire [31:0] dataInProc75West;

	 //Processor 75 control and data signals
	wire wrProc75West;
	wire fullProc75West;
	wire [31:0] dataOutProc75West;

	//Processor 76 control and data signals
	wire rdProc76North;
	wire emptyProc76North;
	wire [31:0] dataInProc76North;

	 //Processor 76 control and data signals
	wire wrProc76North;
	wire fullProc76North;
	wire [31:0] dataOutProc76North;

	 //Processor 76 control and data signals
	wire rdProc76South;
	wire emptyProc76South;
	wire [31:0] dataInProc76South;
	
	 //Processor 76 control and data signals
	wire wrProc76South;
	wire fullProc76South;
	wire [31:0] dataOutProc76South;

	 //Processor 76 control and data signals
	wire rdProc76East;
	wire emptyProc76East;
	wire [31:0] dataInProc76East;
	
	 //Processor 76 control and data signals
	wire wrProc76East;
	wire fullProc76East;
	wire [31:0] dataOutProc76East;

	 //Processor 76 control and data signals
	wire rdProc76West;
	wire emptyProc76West;
	wire [31:0] dataInProc76West;

	 //Processor 76 control and data signals
	wire wrProc76West;
	wire fullProc76West;
	wire [31:0] dataOutProc76West;

	//Processor 77 control and data signals
	wire wrProc77North;
	wire fullProc77North;
	wire [31:0] dataOutProc77North;

	//Processor 77 control and data signals
        wire rdProc77North;
        wire emptyProc77North;
        wire [31:0] dataInProc77North;

	//Processor 77 control and data signals
	wire rdProc77South;
	wire emptyProc77South;
	wire [31:0] dataInProc77South;
		
	 //Processor 77 control and data signals
	wire wrProc77South;
	wire fullProc77South;
	wire [31:0] dataOutProc77South;

	 //Processor 77 control and data signals
	wire wrProc77West;
	wire fullProc77West;
	wire [31:0] dataOutProc77West;
	
	 //Processor 77 control and data signals
	wire rdProc77West;
	wire emptyProc77West;
	wire [31:0] dataInProc77West;

	//Processor 78 control and data signals
	wire wrProc78North;
	wire fullProc78North;
	wire [31:0] dataOutProc78North;

	 //Processor 78 control and data signals
	wire rdProc78North;
	wire emptyProc78North;
	wire [31:0] dataInProc78North;
	
	 //Processor 78 control and data signals
	wire rdProc78South;
	wire emptyProc78South;
	wire [31:0] dataInProc78South;
	
	 //Processor 78 control and data signals
	wire wrProc78South;
	wire fullProc78South;
	wire [31:0] dataOutProc78South;
	
	 //Processor 78 control and data signals
	wire rdProc78East;
	wire emptyProc78East;
	wire [31:0] dataInProc78East;

	 //Processor 78 control and data signals
	wire wrProc78East;
	wire fullProc78East;
	wire [31:0] dataOutProc78East;

	//Processor 79 control and data signals
	wire rdProc79North;
	wire emptyProc79North;
	wire [31:0] dataInProc79North;

	 //Processor 79 control and data signals
	wire wrProc79North;
	wire fullProc79North;
	wire [31:0] dataOutProc79North;

	 //Processor 79 control and data signals
	wire rdProc79South;
	wire emptyProc79South;
	wire [31:0] dataInProc79South;
	
	 //Processor 79 control and data signals
	wire wrProc79South;
	wire fullProc79South;
	wire [31:0] dataOutProc79South;

	 //Processor 79 control and data signals
	wire rdProc79East;
	wire emptyProc79East;
	wire [31:0] dataInProc79East;
	
	 //Processor 79 control and data signals
	wire wrProc79East;
	wire fullProc79East;
	wire [31:0] dataOutProc79East;

	 //Processor 79 control and data signals
	wire rdProc79West;
	wire emptyProc79West;
	wire [31:0] dataInProc79West;

	 //Processor 79 control and data signals
	wire wrProc79West;
	wire fullProc79West;
	wire [31:0] dataOutProc79West;

	//Processor 80 control and data signals
	wire rdProc80North;
	wire emptyProc80North;
	wire [31:0] dataInProc80North;

	 //Processor 80 control and data signals
	wire wrProc80North;
	wire fullProc80North;
	wire [31:0] dataOutProc80North;

	 //Processor 80 control and data signals
	wire rdProc80South;
	wire emptyProc80South;
	wire [31:0] dataInProc80South;
	
	 //Processor 80 control and data signals
	wire wrProc80South;
	wire fullProc80South;
	wire [31:0] dataOutProc80South;

	 //Processor 80 control and data signals
	wire rdProc80East;
	wire emptyProc80East;
	wire [31:0] dataInProc80East;
	
	 //Processor 80 control and data signals
	wire wrProc80East;
	wire fullProc80East;
	wire [31:0] dataOutProc80East;

	 //Processor 80 control and data signals
	wire rdProc80West;
	wire emptyProc80West;
	wire [31:0] dataInProc80West;

	 //Processor 80 control and data signals
	wire wrProc80West;
	wire fullProc80West;
	wire [31:0] dataOutProc80West;

	//Processor 81 control and data signals
	wire rdProc81North;
	wire emptyProc81North;
	wire [31:0] dataInProc81North;

	 //Processor 81 control and data signals
	wire wrProc81North;
	wire fullProc81North;
	wire [31:0] dataOutProc81North;

	 //Processor 81 control and data signals
	wire rdProc81South;
	wire emptyProc81South;
	wire [31:0] dataInProc81South;
	
	 //Processor 81 control and data signals
	wire wrProc81South;
	wire fullProc81South;
	wire [31:0] dataOutProc81South;

	 //Processor 81 control and data signals
	wire rdProc81East;
	wire emptyProc81East;
	wire [31:0] dataInProc81East;
	
	 //Processor 81 control and data signals
	wire wrProc81East;
	wire fullProc81East;
	wire [31:0] dataOutProc81East;

	 //Processor 81 control and data signals
	wire rdProc81West;
	wire emptyProc81West;
	wire [31:0] dataInProc81West;

	 //Processor 81 control and data signals
	wire wrProc81West;
	wire fullProc81West;
	wire [31:0] dataOutProc81West;

	//Processor 82 control and data signals
	wire rdProc82North;
	wire emptyProc82North;
	wire [31:0] dataInProc82North;

	 //Processor 82 control and data signals
	wire wrProc82North;
	wire fullProc82North;
	wire [31:0] dataOutProc82North;

	 //Processor 82 control and data signals
	wire rdProc82South;
	wire emptyProc82South;
	wire [31:0] dataInProc82South;
	
	 //Processor 82 control and data signals
	wire wrProc82South;
	wire fullProc82South;
	wire [31:0] dataOutProc82South;

	 //Processor 82 control and data signals
	wire rdProc82East;
	wire emptyProc82East;
	wire [31:0] dataInProc82East;
	
	 //Processor 82 control and data signals
	wire wrProc82East;
	wire fullProc82East;
	wire [31:0] dataOutProc82East;

	 //Processor 82 control and data signals
	wire rdProc82West;
	wire emptyProc82West;
	wire [31:0] dataInProc82West;

	 //Processor 82 control and data signals
	wire wrProc82West;
	wire fullProc82West;
	wire [31:0] dataOutProc82West;

	//Processor 83 control and data signals
	wire rdProc83North;
	wire emptyProc83North;
	wire [31:0] dataInProc83North;

	 //Processor 83 control and data signals
	wire wrProc83North;
	wire fullProc83North;
	wire [31:0] dataOutProc83North;

	 //Processor 83 control and data signals
	wire rdProc83South;
	wire emptyProc83South;
	wire [31:0] dataInProc83South;
	
	 //Processor 83 control and data signals
	wire wrProc83South;
	wire fullProc83South;
	wire [31:0] dataOutProc83South;

	 //Processor 83 control and data signals
	wire rdProc83East;
	wire emptyProc83East;
	wire [31:0] dataInProc83East;
	
	 //Processor 83 control and data signals
	wire wrProc83East;
	wire fullProc83East;
	wire [31:0] dataOutProc83East;

	 //Processor 83 control and data signals
	wire rdProc83West;
	wire emptyProc83West;
	wire [31:0] dataInProc83West;

	 //Processor 83 control and data signals
	wire wrProc83West;
	wire fullProc83West;
	wire [31:0] dataOutProc83West;

	//Processor 84 control and data signals
	wire rdProc84North;
	wire emptyProc84North;
	wire [31:0] dataInProc84North;

	 //Processor 84 control and data signals
	wire wrProc84North;
	wire fullProc84North;
	wire [31:0] dataOutProc84North;

	 //Processor 84 control and data signals
	wire rdProc84South;
	wire emptyProc84South;
	wire [31:0] dataInProc84South;
	
	 //Processor 84 control and data signals
	wire wrProc84South;
	wire fullProc84South;
	wire [31:0] dataOutProc84South;

	 //Processor 84 control and data signals
	wire rdProc84East;
	wire emptyProc84East;
	wire [31:0] dataInProc84East;
	
	 //Processor 84 control and data signals
	wire wrProc84East;
	wire fullProc84East;
	wire [31:0] dataOutProc84East;

	 //Processor 84 control and data signals
	wire rdProc84West;
	wire emptyProc84West;
	wire [31:0] dataInProc84West;

	 //Processor 84 control and data signals
	wire wrProc84West;
	wire fullProc84West;
	wire [31:0] dataOutProc84West;

	//Processor 85 control and data signals
	wire rdProc85North;
	wire emptyProc85North;
	wire [31:0] dataInProc85North;

	 //Processor 85 control and data signals
	wire wrProc85North;
	wire fullProc85North;
	wire [31:0] dataOutProc85North;

	 //Processor 85 control and data signals
	wire rdProc85South;
	wire emptyProc85South;
	wire [31:0] dataInProc85South;
	
	 //Processor 85 control and data signals
	wire wrProc85South;
	wire fullProc85South;
	wire [31:0] dataOutProc85South;

	 //Processor 85 control and data signals
	wire rdProc85East;
	wire emptyProc85East;
	wire [31:0] dataInProc85East;
	
	 //Processor 85 control and data signals
	wire wrProc85East;
	wire fullProc85East;
	wire [31:0] dataOutProc85East;

	 //Processor 85 control and data signals
	wire rdProc85West;
	wire emptyProc85West;
	wire [31:0] dataInProc85West;

	 //Processor 85 control and data signals
	wire wrProc85West;
	wire fullProc85West;
	wire [31:0] dataOutProc85West;

	//Processor 86 control and data signals
	wire rdProc86North;
	wire emptyProc86North;
	wire [31:0] dataInProc86North;

	 //Processor 86 control and data signals
	wire wrProc86North;
	wire fullProc86North;
	wire [31:0] dataOutProc86North;

	 //Processor 86 control and data signals
	wire rdProc86South;
	wire emptyProc86South;
	wire [31:0] dataInProc86South;
	
	 //Processor 86 control and data signals
	wire wrProc86South;
	wire fullProc86South;
	wire [31:0] dataOutProc86South;

	 //Processor 86 control and data signals
	wire rdProc86East;
	wire emptyProc86East;
	wire [31:0] dataInProc86East;
	
	 //Processor 86 control and data signals
	wire wrProc86East;
	wire fullProc86East;
	wire [31:0] dataOutProc86East;

	 //Processor 86 control and data signals
	wire rdProc86West;
	wire emptyProc86West;
	wire [31:0] dataInProc86West;

	 //Processor 86 control and data signals
	wire wrProc86West;
	wire fullProc86West;
	wire [31:0] dataOutProc86West;

	//Processor 87 control and data signals
	wire rdProc87North;
	wire emptyProc87North;
	wire [31:0] dataInProc87North;

	 //Processor 87 control and data signals
	wire wrProc87North;
	wire fullProc87North;
	wire [31:0] dataOutProc87North;

	 //Processor 87 control and data signals
	wire rdProc87South;
	wire emptyProc87South;
	wire [31:0] dataInProc87South;
	
	 //Processor 87 control and data signals
	wire wrProc87South;
	wire fullProc87South;
	wire [31:0] dataOutProc87South;

	 //Processor 87 control and data signals
	wire rdProc87East;
	wire emptyProc87East;
	wire [31:0] dataInProc87East;
	
	 //Processor 87 control and data signals
	wire wrProc87East;
	wire fullProc87East;
	wire [31:0] dataOutProc87East;

	 //Processor 87 control and data signals
	wire rdProc87West;
	wire emptyProc87West;
	wire [31:0] dataInProc87West;

	 //Processor 87 control and data signals
	wire wrProc87West;
	wire fullProc87West;
	wire [31:0] dataOutProc87West;

	//Processor 88 control and data signals
	wire rdProc88North;
	wire emptyProc88North;
	wire [31:0] dataInProc88North;

	 //Processor 88 control and data signals
	wire wrProc88North;
	wire fullProc88North;
	wire [31:0] dataOutProc88North;

	 //Processor 88 control and data signals
	wire rdProc88South;
	wire emptyProc88South;
	wire [31:0] dataInProc88South;
	
	 //Processor 88 control and data signals
	wire wrProc88South;
	wire fullProc88South;
	wire [31:0] dataOutProc88South;

	 //Processor 88 control and data signals
	wire rdProc88East;
	wire emptyProc88East;
	wire [31:0] dataInProc88East;
	
	 //Processor 88 control and data signals
	wire wrProc88East;
	wire fullProc88East;
	wire [31:0] dataOutProc88East;

	 //Processor 88 control and data signals
	wire rdProc88West;
	wire emptyProc88West;
	wire [31:0] dataInProc88West;

	 //Processor 88 control and data signals
	wire wrProc88West;
	wire fullProc88West;
	wire [31:0] dataOutProc88West;

	//Processor 89 control and data signals
	wire rdProc89North;
	wire emptyProc89North;
	wire [31:0] dataInProc89North;

	 //Processor 89 control and data signals
	wire wrProc89North;
	wire fullProc89North;
	wire [31:0] dataOutProc89North;

	 //Processor 89 control and data signals
	wire rdProc89South;
	wire emptyProc89South;
	wire [31:0] dataInProc89South;
	
	 //Processor 89 control and data signals
	wire wrProc89South;
	wire fullProc89South;
	wire [31:0] dataOutProc89South;

	 //Processor 89 control and data signals
	wire rdProc89East;
	wire emptyProc89East;
	wire [31:0] dataInProc89East;
	
	 //Processor 89 control and data signals
	wire wrProc89East;
	wire fullProc89East;
	wire [31:0] dataOutProc89East;

	 //Processor 89 control and data signals
	wire rdProc89West;
	wire emptyProc89West;
	wire [31:0] dataInProc89West;

	 //Processor 89 control and data signals
	wire wrProc89West;
	wire fullProc89West;
	wire [31:0] dataOutProc89West;

	//Processor 90 control and data signals
	wire wrProc90North;
	wire fullProc90North;
	wire [31:0] dataOutProc90North;

	//Processor 90 control and data signals
        wire rdProc90North;
        wire emptyProc90North;
        wire [31:0] dataInProc90North;

	//Processor 90 control and data signals
	wire rdProc90South;
	wire emptyProc90South;
	wire [31:0] dataInProc90South;
		
	 //Processor 90 control and data signals
	wire wrProc90South;
	wire fullProc90South;
	wire [31:0] dataOutProc90South;

	 //Processor 90 control and data signals
	wire wrProc90West;
	wire fullProc90West;
	wire [31:0] dataOutProc90West;
	
	 //Processor 90 control and data signals
	wire rdProc90West;
	wire emptyProc90West;
	wire [31:0] dataInProc90West;

	//Processor 91 control and data signals
	wire wrProc91North;
	wire fullProc91North;
	wire [31:0] dataOutProc91North;

	 //Processor 91 control and data signals
	wire rdProc91North;
	wire emptyProc91North;
	wire [31:0] dataInProc91North;
	
	 //Processor 91 control and data signals
	wire rdProc91South;
	wire emptyProc91South;
	wire [31:0] dataInProc91South;
	
	 //Processor 91 control and data signals
	wire wrProc91South;
	wire fullProc91South;
	wire [31:0] dataOutProc91South;
	
	 //Processor 91 control and data signals
	wire rdProc91East;
	wire emptyProc91East;
	wire [31:0] dataInProc91East;

	 //Processor 91 control and data signals
	wire wrProc91East;
	wire fullProc91East;
	wire [31:0] dataOutProc91East;

	//Processor 92 control and data signals
	wire rdProc92North;
	wire emptyProc92North;
	wire [31:0] dataInProc92North;

	 //Processor 92 control and data signals
	wire wrProc92North;
	wire fullProc92North;
	wire [31:0] dataOutProc92North;

	 //Processor 92 control and data signals
	wire rdProc92South;
	wire emptyProc92South;
	wire [31:0] dataInProc92South;
	
	 //Processor 92 control and data signals
	wire wrProc92South;
	wire fullProc92South;
	wire [31:0] dataOutProc92South;

	 //Processor 92 control and data signals
	wire rdProc92East;
	wire emptyProc92East;
	wire [31:0] dataInProc92East;
	
	 //Processor 92 control and data signals
	wire wrProc92East;
	wire fullProc92East;
	wire [31:0] dataOutProc92East;

	 //Processor 92 control and data signals
	wire rdProc92West;
	wire emptyProc92West;
	wire [31:0] dataInProc92West;

	 //Processor 92 control and data signals
	wire wrProc92West;
	wire fullProc92West;
	wire [31:0] dataOutProc92West;

	//Processor 93 control and data signals
	wire rdProc93North;
	wire emptyProc93North;
	wire [31:0] dataInProc93North;

	 //Processor 93 control and data signals
	wire wrProc93North;
	wire fullProc93North;
	wire [31:0] dataOutProc93North;

	 //Processor 93 control and data signals
	wire rdProc93South;
	wire emptyProc93South;
	wire [31:0] dataInProc93South;
	
	 //Processor 93 control and data signals
	wire wrProc93South;
	wire fullProc93South;
	wire [31:0] dataOutProc93South;

	 //Processor 93 control and data signals
	wire rdProc93East;
	wire emptyProc93East;
	wire [31:0] dataInProc93East;
	
	 //Processor 93 control and data signals
	wire wrProc93East;
	wire fullProc93East;
	wire [31:0] dataOutProc93East;

	 //Processor 93 control and data signals
	wire rdProc93West;
	wire emptyProc93West;
	wire [31:0] dataInProc93West;

	 //Processor 93 control and data signals
	wire wrProc93West;
	wire fullProc93West;
	wire [31:0] dataOutProc93West;

	//Processor 94 control and data signals
	wire rdProc94North;
	wire emptyProc94North;
	wire [31:0] dataInProc94North;

	 //Processor 94 control and data signals
	wire wrProc94North;
	wire fullProc94North;
	wire [31:0] dataOutProc94North;

	 //Processor 94 control and data signals
	wire rdProc94South;
	wire emptyProc94South;
	wire [31:0] dataInProc94South;
	
	 //Processor 94 control and data signals
	wire wrProc94South;
	wire fullProc94South;
	wire [31:0] dataOutProc94South;

	 //Processor 94 control and data signals
	wire rdProc94East;
	wire emptyProc94East;
	wire [31:0] dataInProc94East;
	
	 //Processor 94 control and data signals
	wire wrProc94East;
	wire fullProc94East;
	wire [31:0] dataOutProc94East;

	 //Processor 94 control and data signals
	wire rdProc94West;
	wire emptyProc94West;
	wire [31:0] dataInProc94West;

	 //Processor 94 control and data signals
	wire wrProc94West;
	wire fullProc94West;
	wire [31:0] dataOutProc94West;

	//Processor 95 control and data signals
	wire rdProc95North;
	wire emptyProc95North;
	wire [31:0] dataInProc95North;

	 //Processor 95 control and data signals
	wire wrProc95North;
	wire fullProc95North;
	wire [31:0] dataOutProc95North;

	 //Processor 95 control and data signals
	wire rdProc95South;
	wire emptyProc95South;
	wire [31:0] dataInProc95South;
	
	 //Processor 95 control and data signals
	wire wrProc95South;
	wire fullProc95South;
	wire [31:0] dataOutProc95South;

	 //Processor 95 control and data signals
	wire rdProc95East;
	wire emptyProc95East;
	wire [31:0] dataInProc95East;
	
	 //Processor 95 control and data signals
	wire wrProc95East;
	wire fullProc95East;
	wire [31:0] dataOutProc95East;

	 //Processor 95 control and data signals
	wire rdProc95West;
	wire emptyProc95West;
	wire [31:0] dataInProc95West;

	 //Processor 95 control and data signals
	wire wrProc95West;
	wire fullProc95West;
	wire [31:0] dataOutProc95West;

	//Processor 96 control and data signals
	wire rdProc96North;
	wire emptyProc96North;
	wire [31:0] dataInProc96North;

	 //Processor 96 control and data signals
	wire wrProc96North;
	wire fullProc96North;
	wire [31:0] dataOutProc96North;

	 //Processor 96 control and data signals
	wire rdProc96South;
	wire emptyProc96South;
	wire [31:0] dataInProc96South;
	
	 //Processor 96 control and data signals
	wire wrProc96South;
	wire fullProc96South;
	wire [31:0] dataOutProc96South;

	 //Processor 96 control and data signals
	wire rdProc96East;
	wire emptyProc96East;
	wire [31:0] dataInProc96East;
	
	 //Processor 96 control and data signals
	wire wrProc96East;
	wire fullProc96East;
	wire [31:0] dataOutProc96East;

	 //Processor 96 control and data signals
	wire rdProc96West;
	wire emptyProc96West;
	wire [31:0] dataInProc96West;

	 //Processor 96 control and data signals
	wire wrProc96West;
	wire fullProc96West;
	wire [31:0] dataOutProc96West;

	//Processor 97 control and data signals
	wire rdProc97North;
	wire emptyProc97North;
	wire [31:0] dataInProc97North;

	 //Processor 97 control and data signals
	wire wrProc97North;
	wire fullProc97North;
	wire [31:0] dataOutProc97North;

	 //Processor 97 control and data signals
	wire rdProc97South;
	wire emptyProc97South;
	wire [31:0] dataInProc97South;
	
	 //Processor 97 control and data signals
	wire wrProc97South;
	wire fullProc97South;
	wire [31:0] dataOutProc97South;

	 //Processor 97 control and data signals
	wire rdProc97East;
	wire emptyProc97East;
	wire [31:0] dataInProc97East;
	
	 //Processor 97 control and data signals
	wire wrProc97East;
	wire fullProc97East;
	wire [31:0] dataOutProc97East;

	 //Processor 97 control and data signals
	wire rdProc97West;
	wire emptyProc97West;
	wire [31:0] dataInProc97West;

	 //Processor 97 control and data signals
	wire wrProc97West;
	wire fullProc97West;
	wire [31:0] dataOutProc97West;

	//Processor 98 control and data signals
	wire rdProc98North;
	wire emptyProc98North;
	wire [31:0] dataInProc98North;

	 //Processor 98 control and data signals
	wire wrProc98North;
	wire fullProc98North;
	wire [31:0] dataOutProc98North;

	 //Processor 98 control and data signals
	wire rdProc98South;
	wire emptyProc98South;
	wire [31:0] dataInProc98South;
	
	 //Processor 98 control and data signals
	wire wrProc98South;
	wire fullProc98South;
	wire [31:0] dataOutProc98South;

	 //Processor 98 control and data signals
	wire rdProc98East;
	wire emptyProc98East;
	wire [31:0] dataInProc98East;
	
	 //Processor 98 control and data signals
	wire wrProc98East;
	wire fullProc98East;
	wire [31:0] dataOutProc98East;

	 //Processor 98 control and data signals
	wire rdProc98West;
	wire emptyProc98West;
	wire [31:0] dataInProc98West;

	 //Processor 98 control and data signals
	wire wrProc98West;
	wire fullProc98West;
	wire [31:0] dataOutProc98West;

	//Processor 99 control and data signals
	wire rdProc99North;
	wire emptyProc99North;
	wire [31:0] dataInProc99North;

	 //Processor 99 control and data signals
	wire wrProc99North;
	wire fullProc99North;
	wire [31:0] dataOutProc99North;

	 //Processor 99 control and data signals
	wire rdProc99South;
	wire emptyProc99South;
	wire [31:0] dataInProc99South;
	
	 //Processor 99 control and data signals
	wire wrProc99South;
	wire fullProc99South;
	wire [31:0] dataOutProc99South;

	 //Processor 99 control and data signals
	wire rdProc99East;
	wire emptyProc99East;
	wire [31:0] dataInProc99East;
	
	 //Processor 99 control and data signals
	wire wrProc99East;
	wire fullProc99East;
	wire [31:0] dataOutProc99East;

	 //Processor 99 control and data signals
	wire rdProc99West;
	wire emptyProc99West;
	wire [31:0] dataInProc99West;

	 //Processor 99 control and data signals
	wire wrProc99West;
	wire fullProc99West;
	wire [31:0] dataOutProc99West;

	//Processor 100 control and data signals
	wire rdProc100North;
	wire emptyProc100North;
	wire [31:0] dataInProc100North;

	 //Processor 100 control and data signals
	wire wrProc100North;
	wire fullProc100North;
	wire [31:0] dataOutProc100North;

	 //Processor 100 control and data signals
	wire rdProc100South;
	wire emptyProc100South;
	wire [31:0] dataInProc100South;
	
	 //Processor 100 control and data signals
	wire wrProc100South;
	wire fullProc100South;
	wire [31:0] dataOutProc100South;

	 //Processor 100 control and data signals
	wire rdProc100East;
	wire emptyProc100East;
	wire [31:0] dataInProc100East;
	
	 //Processor 100 control and data signals
	wire wrProc100East;
	wire fullProc100East;
	wire [31:0] dataOutProc100East;

	 //Processor 100 control and data signals
	wire rdProc100West;
	wire emptyProc100West;
	wire [31:0] dataInProc100West;

	 //Processor 100 control and data signals
	wire wrProc100West;
	wire fullProc100West;
	wire [31:0] dataOutProc100West;

	//Processor 101 control and data signals
	wire rdProc101North;
	wire emptyProc101North;
	wire [31:0] dataInProc101North;

	 //Processor 101 control and data signals
	wire wrProc101North;
	wire fullProc101North;
	wire [31:0] dataOutProc101North;

	 //Processor 101 control and data signals
	wire rdProc101South;
	wire emptyProc101South;
	wire [31:0] dataInProc101South;
	
	 //Processor 101 control and data signals
	wire wrProc101South;
	wire fullProc101South;
	wire [31:0] dataOutProc101South;

	 //Processor 101 control and data signals
	wire rdProc101East;
	wire emptyProc101East;
	wire [31:0] dataInProc101East;
	
	 //Processor 101 control and data signals
	wire wrProc101East;
	wire fullProc101East;
	wire [31:0] dataOutProc101East;

	 //Processor 101 control and data signals
	wire rdProc101West;
	wire emptyProc101West;
	wire [31:0] dataInProc101West;

	 //Processor 101 control and data signals
	wire wrProc101West;
	wire fullProc101West;
	wire [31:0] dataOutProc101West;

	//Processor 102 control and data signals
	wire rdProc102North;
	wire emptyProc102North;
	wire [31:0] dataInProc102North;

	 //Processor 102 control and data signals
	wire wrProc102North;
	wire fullProc102North;
	wire [31:0] dataOutProc102North;

	 //Processor 102 control and data signals
	wire rdProc102South;
	wire emptyProc102South;
	wire [31:0] dataInProc102South;
	
	 //Processor 102 control and data signals
	wire wrProc102South;
	wire fullProc102South;
	wire [31:0] dataOutProc102South;

	 //Processor 102 control and data signals
	wire rdProc102East;
	wire emptyProc102East;
	wire [31:0] dataInProc102East;
	
	 //Processor 102 control and data signals
	wire wrProc102East;
	wire fullProc102East;
	wire [31:0] dataOutProc102East;

	 //Processor 102 control and data signals
	wire rdProc102West;
	wire emptyProc102West;
	wire [31:0] dataInProc102West;

	 //Processor 102 control and data signals
	wire wrProc102West;
	wire fullProc102West;
	wire [31:0] dataOutProc102West;

	//Processor 103 control and data signals
	wire wrProc103North;
	wire fullProc103North;
	wire [31:0] dataOutProc103North;

	//Processor 103 control and data signals
        wire rdProc103North;
        wire emptyProc103North;
        wire [31:0] dataInProc103North;

	//Processor 103 control and data signals
	wire rdProc103South;
	wire emptyProc103South;
	wire [31:0] dataInProc103South;
		
	 //Processor 103 control and data signals
	wire wrProc103South;
	wire fullProc103South;
	wire [31:0] dataOutProc103South;

	 //Processor 103 control and data signals
	wire wrProc103West;
	wire fullProc103West;
	wire [31:0] dataOutProc103West;
	
	 //Processor 103 control and data signals
	wire rdProc103West;
	wire emptyProc103West;
	wire [31:0] dataInProc103West;

	//Processor 104 control and data signals
	wire wrProc104North;
	wire fullProc104North;
	wire [31:0] dataOutProc104North;

	 //Processor 104 control and data signals
	wire rdProc104North;
	wire emptyProc104North;
	wire [31:0] dataInProc104North;
	
	 //Processor 104 control and data signals
	wire rdProc104South;
	wire emptyProc104South;
	wire [31:0] dataInProc104South;
	
	 //Processor 104 control and data signals
	wire wrProc104South;
	wire fullProc104South;
	wire [31:0] dataOutProc104South;
	
	 //Processor 104 control and data signals
	wire rdProc104East;
	wire emptyProc104East;
	wire [31:0] dataInProc104East;

	 //Processor 104 control and data signals
	wire wrProc104East;
	wire fullProc104East;
	wire [31:0] dataOutProc104East;

	//Processor 105 control and data signals
	wire rdProc105North;
	wire emptyProc105North;
	wire [31:0] dataInProc105North;

	 //Processor 105 control and data signals
	wire wrProc105North;
	wire fullProc105North;
	wire [31:0] dataOutProc105North;

	 //Processor 105 control and data signals
	wire rdProc105South;
	wire emptyProc105South;
	wire [31:0] dataInProc105South;
	
	 //Processor 105 control and data signals
	wire wrProc105South;
	wire fullProc105South;
	wire [31:0] dataOutProc105South;

	 //Processor 105 control and data signals
	wire rdProc105East;
	wire emptyProc105East;
	wire [31:0] dataInProc105East;
	
	 //Processor 105 control and data signals
	wire wrProc105East;
	wire fullProc105East;
	wire [31:0] dataOutProc105East;

	 //Processor 105 control and data signals
	wire rdProc105West;
	wire emptyProc105West;
	wire [31:0] dataInProc105West;

	 //Processor 105 control and data signals
	wire wrProc105West;
	wire fullProc105West;
	wire [31:0] dataOutProc105West;

	//Processor 106 control and data signals
	wire rdProc106North;
	wire emptyProc106North;
	wire [31:0] dataInProc106North;

	 //Processor 106 control and data signals
	wire wrProc106North;
	wire fullProc106North;
	wire [31:0] dataOutProc106North;

	 //Processor 106 control and data signals
	wire rdProc106South;
	wire emptyProc106South;
	wire [31:0] dataInProc106South;
	
	 //Processor 106 control and data signals
	wire wrProc106South;
	wire fullProc106South;
	wire [31:0] dataOutProc106South;

	 //Processor 106 control and data signals
	wire rdProc106East;
	wire emptyProc106East;
	wire [31:0] dataInProc106East;
	
	 //Processor 106 control and data signals
	wire wrProc106East;
	wire fullProc106East;
	wire [31:0] dataOutProc106East;

	 //Processor 106 control and data signals
	wire rdProc106West;
	wire emptyProc106West;
	wire [31:0] dataInProc106West;

	 //Processor 106 control and data signals
	wire wrProc106West;
	wire fullProc106West;
	wire [31:0] dataOutProc106West;

	//Processor 107 control and data signals
	wire rdProc107North;
	wire emptyProc107North;
	wire [31:0] dataInProc107North;

	 //Processor 107 control and data signals
	wire wrProc107North;
	wire fullProc107North;
	wire [31:0] dataOutProc107North;

	 //Processor 107 control and data signals
	wire rdProc107South;
	wire emptyProc107South;
	wire [31:0] dataInProc107South;
	
	 //Processor 107 control and data signals
	wire wrProc107South;
	wire fullProc107South;
	wire [31:0] dataOutProc107South;

	 //Processor 107 control and data signals
	wire rdProc107East;
	wire emptyProc107East;
	wire [31:0] dataInProc107East;
	
	 //Processor 107 control and data signals
	wire wrProc107East;
	wire fullProc107East;
	wire [31:0] dataOutProc107East;

	 //Processor 107 control and data signals
	wire rdProc107West;
	wire emptyProc107West;
	wire [31:0] dataInProc107West;

	 //Processor 107 control and data signals
	wire wrProc107West;
	wire fullProc107West;
	wire [31:0] dataOutProc107West;

	//Processor 108 control and data signals
	wire rdProc108North;
	wire emptyProc108North;
	wire [31:0] dataInProc108North;

	 //Processor 108 control and data signals
	wire wrProc108North;
	wire fullProc108North;
	wire [31:0] dataOutProc108North;

	 //Processor 108 control and data signals
	wire rdProc108South;
	wire emptyProc108South;
	wire [31:0] dataInProc108South;
	
	 //Processor 108 control and data signals
	wire wrProc108South;
	wire fullProc108South;
	wire [31:0] dataOutProc108South;

	 //Processor 108 control and data signals
	wire rdProc108East;
	wire emptyProc108East;
	wire [31:0] dataInProc108East;
	
	 //Processor 108 control and data signals
	wire wrProc108East;
	wire fullProc108East;
	wire [31:0] dataOutProc108East;

	 //Processor 108 control and data signals
	wire rdProc108West;
	wire emptyProc108West;
	wire [31:0] dataInProc108West;

	 //Processor 108 control and data signals
	wire wrProc108West;
	wire fullProc108West;
	wire [31:0] dataOutProc108West;

	//Processor 109 control and data signals
	wire rdProc109North;
	wire emptyProc109North;
	wire [31:0] dataInProc109North;

	 //Processor 109 control and data signals
	wire wrProc109North;
	wire fullProc109North;
	wire [31:0] dataOutProc109North;

	 //Processor 109 control and data signals
	wire rdProc109South;
	wire emptyProc109South;
	wire [31:0] dataInProc109South;
	
	 //Processor 109 control and data signals
	wire wrProc109South;
	wire fullProc109South;
	wire [31:0] dataOutProc109South;

	 //Processor 109 control and data signals
	wire rdProc109East;
	wire emptyProc109East;
	wire [31:0] dataInProc109East;
	
	 //Processor 109 control and data signals
	wire wrProc109East;
	wire fullProc109East;
	wire [31:0] dataOutProc109East;

	 //Processor 109 control and data signals
	wire rdProc109West;
	wire emptyProc109West;
	wire [31:0] dataInProc109West;

	 //Processor 109 control and data signals
	wire wrProc109West;
	wire fullProc109West;
	wire [31:0] dataOutProc109West;

	//Processor 110 control and data signals
	wire rdProc110North;
	wire emptyProc110North;
	wire [31:0] dataInProc110North;

	 //Processor 110 control and data signals
	wire wrProc110North;
	wire fullProc110North;
	wire [31:0] dataOutProc110North;

	 //Processor 110 control and data signals
	wire rdProc110South;
	wire emptyProc110South;
	wire [31:0] dataInProc110South;
	
	 //Processor 110 control and data signals
	wire wrProc110South;
	wire fullProc110South;
	wire [31:0] dataOutProc110South;

	 //Processor 110 control and data signals
	wire rdProc110East;
	wire emptyProc110East;
	wire [31:0] dataInProc110East;
	
	 //Processor 110 control and data signals
	wire wrProc110East;
	wire fullProc110East;
	wire [31:0] dataOutProc110East;

	 //Processor 110 control and data signals
	wire rdProc110West;
	wire emptyProc110West;
	wire [31:0] dataInProc110West;

	 //Processor 110 control and data signals
	wire wrProc110West;
	wire fullProc110West;
	wire [31:0] dataOutProc110West;

	//Processor 111 control and data signals
	wire rdProc111North;
	wire emptyProc111North;
	wire [31:0] dataInProc111North;

	 //Processor 111 control and data signals
	wire wrProc111North;
	wire fullProc111North;
	wire [31:0] dataOutProc111North;

	 //Processor 111 control and data signals
	wire rdProc111South;
	wire emptyProc111South;
	wire [31:0] dataInProc111South;
	
	 //Processor 111 control and data signals
	wire wrProc111South;
	wire fullProc111South;
	wire [31:0] dataOutProc111South;

	 //Processor 111 control and data signals
	wire rdProc111East;
	wire emptyProc111East;
	wire [31:0] dataInProc111East;
	
	 //Processor 111 control and data signals
	wire wrProc111East;
	wire fullProc111East;
	wire [31:0] dataOutProc111East;

	 //Processor 111 control and data signals
	wire rdProc111West;
	wire emptyProc111West;
	wire [31:0] dataInProc111West;

	 //Processor 111 control and data signals
	wire wrProc111West;
	wire fullProc111West;
	wire [31:0] dataOutProc111West;

	//Processor 112 control and data signals
	wire rdProc112North;
	wire emptyProc112North;
	wire [31:0] dataInProc112North;

	 //Processor 112 control and data signals
	wire wrProc112North;
	wire fullProc112North;
	wire [31:0] dataOutProc112North;

	 //Processor 112 control and data signals
	wire rdProc112South;
	wire emptyProc112South;
	wire [31:0] dataInProc112South;
	
	 //Processor 112 control and data signals
	wire wrProc112South;
	wire fullProc112South;
	wire [31:0] dataOutProc112South;

	 //Processor 112 control and data signals
	wire rdProc112East;
	wire emptyProc112East;
	wire [31:0] dataInProc112East;
	
	 //Processor 112 control and data signals
	wire wrProc112East;
	wire fullProc112East;
	wire [31:0] dataOutProc112East;

	 //Processor 112 control and data signals
	wire rdProc112West;
	wire emptyProc112West;
	wire [31:0] dataInProc112West;

	 //Processor 112 control and data signals
	wire wrProc112West;
	wire fullProc112West;
	wire [31:0] dataOutProc112West;

	//Processor 113 control and data signals
	wire rdProc113North;
	wire emptyProc113North;
	wire [31:0] dataInProc113North;

	 //Processor 113 control and data signals
	wire wrProc113North;
	wire fullProc113North;
	wire [31:0] dataOutProc113North;

	 //Processor 113 control and data signals
	wire rdProc113South;
	wire emptyProc113South;
	wire [31:0] dataInProc113South;
	
	 //Processor 113 control and data signals
	wire wrProc113South;
	wire fullProc113South;
	wire [31:0] dataOutProc113South;

	 //Processor 113 control and data signals
	wire rdProc113East;
	wire emptyProc113East;
	wire [31:0] dataInProc113East;
	
	 //Processor 113 control and data signals
	wire wrProc113East;
	wire fullProc113East;
	wire [31:0] dataOutProc113East;

	 //Processor 113 control and data signals
	wire rdProc113West;
	wire emptyProc113West;
	wire [31:0] dataInProc113West;

	 //Processor 113 control and data signals
	wire wrProc113West;
	wire fullProc113West;
	wire [31:0] dataOutProc113West;

	//Processor 114 control and data signals
	wire rdProc114North;
	wire emptyProc114North;
	wire [31:0] dataInProc114North;

	 //Processor 114 control and data signals
	wire wrProc114North;
	wire fullProc114North;
	wire [31:0] dataOutProc114North;

	 //Processor 114 control and data signals
	wire rdProc114South;
	wire emptyProc114South;
	wire [31:0] dataInProc114South;
	
	 //Processor 114 control and data signals
	wire wrProc114South;
	wire fullProc114South;
	wire [31:0] dataOutProc114South;

	 //Processor 114 control and data signals
	wire rdProc114East;
	wire emptyProc114East;
	wire [31:0] dataInProc114East;
	
	 //Processor 114 control and data signals
	wire wrProc114East;
	wire fullProc114East;
	wire [31:0] dataOutProc114East;

	 //Processor 114 control and data signals
	wire rdProc114West;
	wire emptyProc114West;
	wire [31:0] dataInProc114West;

	 //Processor 114 control and data signals
	wire wrProc114West;
	wire fullProc114West;
	wire [31:0] dataOutProc114West;

	//Processor 115 control and data signals
	wire rdProc115North;
	wire emptyProc115North;
	wire [31:0] dataInProc115North;

	 //Processor 115 control and data signals
	wire wrProc115North;
	wire fullProc115North;
	wire [31:0] dataOutProc115North;

	 //Processor 115 control and data signals
	wire rdProc115South;
	wire emptyProc115South;
	wire [31:0] dataInProc115South;
	
	 //Processor 115 control and data signals
	wire wrProc115South;
	wire fullProc115South;
	wire [31:0] dataOutProc115South;

	 //Processor 115 control and data signals
	wire rdProc115East;
	wire emptyProc115East;
	wire [31:0] dataInProc115East;
	
	 //Processor 115 control and data signals
	wire wrProc115East;
	wire fullProc115East;
	wire [31:0] dataOutProc115East;

	 //Processor 115 control and data signals
	wire rdProc115West;
	wire emptyProc115West;
	wire [31:0] dataInProc115West;

	 //Processor 115 control and data signals
	wire wrProc115West;
	wire fullProc115West;
	wire [31:0] dataOutProc115West;

	//Processor 116 control and data signals
	wire wrProc116North;
	wire fullProc116North;
	wire [31:0] dataOutProc116North;

	//Processor 116 control and data signals
        wire rdProc116North;
        wire emptyProc116North;
        wire [31:0] dataInProc116North;

	//Processor 116 control and data signals
	wire rdProc116South;
	wire emptyProc116South;
	wire [31:0] dataInProc116South;
		
	 //Processor 116 control and data signals
	wire wrProc116South;
	wire fullProc116South;
	wire [31:0] dataOutProc116South;

	 //Processor 116 control and data signals
	wire wrProc116West;
	wire fullProc116West;
	wire [31:0] dataOutProc116West;
	
	 //Processor 116 control and data signals
	wire rdProc116West;
	wire emptyProc116West;
	wire [31:0] dataInProc116West;

	//Processor 117 control and data signals
	wire wrProc117North;
	wire fullProc117North;
	wire [31:0] dataOutProc117North;

	 //Processor 117 control and data signals
	wire rdProc117North;
	wire emptyProc117North;
	wire [31:0] dataInProc117North;
	
	 //Processor 117 control and data signals
	wire rdProc117South;
	wire emptyProc117South;
	wire [31:0] dataInProc117South;
	
	 //Processor 117 control and data signals
	wire wrProc117South;
	wire fullProc117South;
	wire [31:0] dataOutProc117South;
	
	 //Processor 117 control and data signals
	wire rdProc117East;
	wire emptyProc117East;
	wire [31:0] dataInProc117East;

	 //Processor 117 control and data signals
	wire wrProc117East;
	wire fullProc117East;
	wire [31:0] dataOutProc117East;

	//Processor 118 control and data signals
	wire rdProc118North;
	wire emptyProc118North;
	wire [31:0] dataInProc118North;

	 //Processor 118 control and data signals
	wire wrProc118North;
	wire fullProc118North;
	wire [31:0] dataOutProc118North;

	 //Processor 118 control and data signals
	wire rdProc118South;
	wire emptyProc118South;
	wire [31:0] dataInProc118South;
	
	 //Processor 118 control and data signals
	wire wrProc118South;
	wire fullProc118South;
	wire [31:0] dataOutProc118South;

	 //Processor 118 control and data signals
	wire rdProc118East;
	wire emptyProc118East;
	wire [31:0] dataInProc118East;
	
	 //Processor 118 control and data signals
	wire wrProc118East;
	wire fullProc118East;
	wire [31:0] dataOutProc118East;

	 //Processor 118 control and data signals
	wire rdProc118West;
	wire emptyProc118West;
	wire [31:0] dataInProc118West;

	 //Processor 118 control and data signals
	wire wrProc118West;
	wire fullProc118West;
	wire [31:0] dataOutProc118West;

	//Processor 119 control and data signals
	wire rdProc119North;
	wire emptyProc119North;
	wire [31:0] dataInProc119North;

	 //Processor 119 control and data signals
	wire wrProc119North;
	wire fullProc119North;
	wire [31:0] dataOutProc119North;

	 //Processor 119 control and data signals
	wire rdProc119South;
	wire emptyProc119South;
	wire [31:0] dataInProc119South;
	
	 //Processor 119 control and data signals
	wire wrProc119South;
	wire fullProc119South;
	wire [31:0] dataOutProc119South;

	 //Processor 119 control and data signals
	wire rdProc119East;
	wire emptyProc119East;
	wire [31:0] dataInProc119East;
	
	 //Processor 119 control and data signals
	wire wrProc119East;
	wire fullProc119East;
	wire [31:0] dataOutProc119East;

	 //Processor 119 control and data signals
	wire rdProc119West;
	wire emptyProc119West;
	wire [31:0] dataInProc119West;

	 //Processor 119 control and data signals
	wire wrProc119West;
	wire fullProc119West;
	wire [31:0] dataOutProc119West;

	//Processor 120 control and data signals
	wire rdProc120North;
	wire emptyProc120North;
	wire [31:0] dataInProc120North;

	 //Processor 120 control and data signals
	wire wrProc120North;
	wire fullProc120North;
	wire [31:0] dataOutProc120North;

	 //Processor 120 control and data signals
	wire rdProc120South;
	wire emptyProc120South;
	wire [31:0] dataInProc120South;
	
	 //Processor 120 control and data signals
	wire wrProc120South;
	wire fullProc120South;
	wire [31:0] dataOutProc120South;

	 //Processor 120 control and data signals
	wire rdProc120East;
	wire emptyProc120East;
	wire [31:0] dataInProc120East;
	
	 //Processor 120 control and data signals
	wire wrProc120East;
	wire fullProc120East;
	wire [31:0] dataOutProc120East;

	 //Processor 120 control and data signals
	wire rdProc120West;
	wire emptyProc120West;
	wire [31:0] dataInProc120West;

	 //Processor 120 control and data signals
	wire wrProc120West;
	wire fullProc120West;
	wire [31:0] dataOutProc120West;

	//Processor 121 control and data signals
	wire rdProc121North;
	wire emptyProc121North;
	wire [31:0] dataInProc121North;

	 //Processor 121 control and data signals
	wire wrProc121North;
	wire fullProc121North;
	wire [31:0] dataOutProc121North;

	 //Processor 121 control and data signals
	wire rdProc121South;
	wire emptyProc121South;
	wire [31:0] dataInProc121South;
	
	 //Processor 121 control and data signals
	wire wrProc121South;
	wire fullProc121South;
	wire [31:0] dataOutProc121South;

	 //Processor 121 control and data signals
	wire rdProc121East;
	wire emptyProc121East;
	wire [31:0] dataInProc121East;
	
	 //Processor 121 control and data signals
	wire wrProc121East;
	wire fullProc121East;
	wire [31:0] dataOutProc121East;

	 //Processor 121 control and data signals
	wire rdProc121West;
	wire emptyProc121West;
	wire [31:0] dataInProc121West;

	 //Processor 121 control and data signals
	wire wrProc121West;
	wire fullProc121West;
	wire [31:0] dataOutProc121West;

	//Processor 122 control and data signals
	wire rdProc122North;
	wire emptyProc122North;
	wire [31:0] dataInProc122North;

	 //Processor 122 control and data signals
	wire wrProc122North;
	wire fullProc122North;
	wire [31:0] dataOutProc122North;

	 //Processor 122 control and data signals
	wire rdProc122South;
	wire emptyProc122South;
	wire [31:0] dataInProc122South;
	
	 //Processor 122 control and data signals
	wire wrProc122South;
	wire fullProc122South;
	wire [31:0] dataOutProc122South;

	 //Processor 122 control and data signals
	wire rdProc122East;
	wire emptyProc122East;
	wire [31:0] dataInProc122East;
	
	 //Processor 122 control and data signals
	wire wrProc122East;
	wire fullProc122East;
	wire [31:0] dataOutProc122East;

	 //Processor 122 control and data signals
	wire rdProc122West;
	wire emptyProc122West;
	wire [31:0] dataInProc122West;

	 //Processor 122 control and data signals
	wire wrProc122West;
	wire fullProc122West;
	wire [31:0] dataOutProc122West;

	//Processor 123 control and data signals
	wire rdProc123North;
	wire emptyProc123North;
	wire [31:0] dataInProc123North;

	 //Processor 123 control and data signals
	wire wrProc123North;
	wire fullProc123North;
	wire [31:0] dataOutProc123North;

	 //Processor 123 control and data signals
	wire rdProc123South;
	wire emptyProc123South;
	wire [31:0] dataInProc123South;
	
	 //Processor 123 control and data signals
	wire wrProc123South;
	wire fullProc123South;
	wire [31:0] dataOutProc123South;

	 //Processor 123 control and data signals
	wire rdProc123East;
	wire emptyProc123East;
	wire [31:0] dataInProc123East;
	
	 //Processor 123 control and data signals
	wire wrProc123East;
	wire fullProc123East;
	wire [31:0] dataOutProc123East;

	 //Processor 123 control and data signals
	wire rdProc123West;
	wire emptyProc123West;
	wire [31:0] dataInProc123West;

	 //Processor 123 control and data signals
	wire wrProc123West;
	wire fullProc123West;
	wire [31:0] dataOutProc123West;

	//Processor 124 control and data signals
	wire rdProc124North;
	wire emptyProc124North;
	wire [31:0] dataInProc124North;

	 //Processor 124 control and data signals
	wire wrProc124North;
	wire fullProc124North;
	wire [31:0] dataOutProc124North;

	 //Processor 124 control and data signals
	wire rdProc124South;
	wire emptyProc124South;
	wire [31:0] dataInProc124South;
	
	 //Processor 124 control and data signals
	wire wrProc124South;
	wire fullProc124South;
	wire [31:0] dataOutProc124South;

	 //Processor 124 control and data signals
	wire rdProc124East;
	wire emptyProc124East;
	wire [31:0] dataInProc124East;
	
	 //Processor 124 control and data signals
	wire wrProc124East;
	wire fullProc124East;
	wire [31:0] dataOutProc124East;

	 //Processor 124 control and data signals
	wire rdProc124West;
	wire emptyProc124West;
	wire [31:0] dataInProc124West;

	 //Processor 124 control and data signals
	wire wrProc124West;
	wire fullProc124West;
	wire [31:0] dataOutProc124West;

	//Processor 125 control and data signals
	wire rdProc125North;
	wire emptyProc125North;
	wire [31:0] dataInProc125North;

	 //Processor 125 control and data signals
	wire wrProc125North;
	wire fullProc125North;
	wire [31:0] dataOutProc125North;

	 //Processor 125 control and data signals
	wire rdProc125South;
	wire emptyProc125South;
	wire [31:0] dataInProc125South;
	
	 //Processor 125 control and data signals
	wire wrProc125South;
	wire fullProc125South;
	wire [31:0] dataOutProc125South;

	 //Processor 125 control and data signals
	wire rdProc125East;
	wire emptyProc125East;
	wire [31:0] dataInProc125East;
	
	 //Processor 125 control and data signals
	wire wrProc125East;
	wire fullProc125East;
	wire [31:0] dataOutProc125East;

	 //Processor 125 control and data signals
	wire rdProc125West;
	wire emptyProc125West;
	wire [31:0] dataInProc125West;

	 //Processor 125 control and data signals
	wire wrProc125West;
	wire fullProc125West;
	wire [31:0] dataOutProc125West;

	//Processor 126 control and data signals
	wire rdProc126North;
	wire emptyProc126North;
	wire [31:0] dataInProc126North;

	 //Processor 126 control and data signals
	wire wrProc126North;
	wire fullProc126North;
	wire [31:0] dataOutProc126North;

	 //Processor 126 control and data signals
	wire rdProc126South;
	wire emptyProc126South;
	wire [31:0] dataInProc126South;
	
	 //Processor 126 control and data signals
	wire wrProc126South;
	wire fullProc126South;
	wire [31:0] dataOutProc126South;

	 //Processor 126 control and data signals
	wire rdProc126East;
	wire emptyProc126East;
	wire [31:0] dataInProc126East;
	
	 //Processor 126 control and data signals
	wire wrProc126East;
	wire fullProc126East;
	wire [31:0] dataOutProc126East;

	 //Processor 126 control and data signals
	wire rdProc126West;
	wire emptyProc126West;
	wire [31:0] dataInProc126West;

	 //Processor 126 control and data signals
	wire wrProc126West;
	wire fullProc126West;
	wire [31:0] dataOutProc126West;

	//Processor 127 control and data signals
	wire rdProc127North;
	wire emptyProc127North;
	wire [31:0] dataInProc127North;

	 //Processor 127 control and data signals
	wire wrProc127North;
	wire fullProc127North;
	wire [31:0] dataOutProc127North;

	 //Processor 127 control and data signals
	wire rdProc127South;
	wire emptyProc127South;
	wire [31:0] dataInProc127South;
	
	 //Processor 127 control and data signals
	wire wrProc127South;
	wire fullProc127South;
	wire [31:0] dataOutProc127South;

	 //Processor 127 control and data signals
	wire rdProc127East;
	wire emptyProc127East;
	wire [31:0] dataInProc127East;
	
	 //Processor 127 control and data signals
	wire wrProc127East;
	wire fullProc127East;
	wire [31:0] dataOutProc127East;

	 //Processor 127 control and data signals
	wire rdProc127West;
	wire emptyProc127West;
	wire [31:0] dataInProc127West;

	 //Processor 127 control and data signals
	wire wrProc127West;
	wire fullProc127West;
	wire [31:0] dataOutProc127West;

	//Processor 128 control and data signals
	wire rdProc128North;
	wire emptyProc128North;
	wire [31:0] dataInProc128North;

	 //Processor 128 control and data signals
	wire wrProc128North;
	wire fullProc128North;
	wire [31:0] dataOutProc128North;

	 //Processor 128 control and data signals
	wire rdProc128South;
	wire emptyProc128South;
	wire [31:0] dataInProc128South;
	
	 //Processor 128 control and data signals
	wire wrProc128South;
	wire fullProc128South;
	wire [31:0] dataOutProc128South;

	 //Processor 128 control and data signals
	wire rdProc128East;
	wire emptyProc128East;
	wire [31:0] dataInProc128East;
	
	 //Processor 128 control and data signals
	wire wrProc128East;
	wire fullProc128East;
	wire [31:0] dataOutProc128East;

	 //Processor 128 control and data signals
	wire rdProc128West;
	wire emptyProc128West;
	wire [31:0] dataInProc128West;

	 //Processor 128 control and data signals
	wire wrProc128West;
	wire fullProc128West;
	wire [31:0] dataOutProc128West;

	//Processor 129 control and data signals
	wire wrProc129North;
	wire fullProc129North;
	wire [31:0] dataOutProc129North;

	//Processor 129 control and data signals
        wire rdProc129North;
        wire emptyProc129North;
        wire [31:0] dataInProc129North;

	//Processor 129 control and data signals
	wire rdProc129South;
	wire emptyProc129South;
	wire [31:0] dataInProc129South;
		
	 //Processor 129 control and data signals
	wire wrProc129South;
	wire fullProc129South;
	wire [31:0] dataOutProc129South;

	 //Processor 129 control and data signals
	wire wrProc129West;
	wire fullProc129West;
	wire [31:0] dataOutProc129West;
	
	 //Processor 129 control and data signals
	wire rdProc129West;
	wire emptyProc129West;
	wire [31:0] dataInProc129West;

	//Processor 130 control and data signals
	wire wrProc130North;
	wire fullProc130North;
	wire [31:0] dataOutProc130North;

	 //Processor 130 control and data signals
	wire rdProc130North;
	wire emptyProc130North;
	wire [31:0] dataInProc130North;
	
	 //Processor 130 control and data signals
	wire rdProc130South;
	wire emptyProc130South;
	wire [31:0] dataInProc130South;
	
	 //Processor 130 control and data signals
	wire wrProc130South;
	wire fullProc130South;
	wire [31:0] dataOutProc130South;
	
	 //Processor 130 control and data signals
	wire rdProc130East;
	wire emptyProc130East;
	wire [31:0] dataInProc130East;

	 //Processor 130 control and data signals
	wire wrProc130East;
	wire fullProc130East;
	wire [31:0] dataOutProc130East;

	//Processor 131 control and data signals
	wire rdProc131North;
	wire emptyProc131North;
	wire [31:0] dataInProc131North;

	 //Processor 131 control and data signals
	wire wrProc131North;
	wire fullProc131North;
	wire [31:0] dataOutProc131North;

	 //Processor 131 control and data signals
	wire rdProc131South;
	wire emptyProc131South;
	wire [31:0] dataInProc131South;
	
	 //Processor 131 control and data signals
	wire wrProc131South;
	wire fullProc131South;
	wire [31:0] dataOutProc131South;

	 //Processor 131 control and data signals
	wire rdProc131East;
	wire emptyProc131East;
	wire [31:0] dataInProc131East;
	
	 //Processor 131 control and data signals
	wire wrProc131East;
	wire fullProc131East;
	wire [31:0] dataOutProc131East;

	 //Processor 131 control and data signals
	wire rdProc131West;
	wire emptyProc131West;
	wire [31:0] dataInProc131West;

	 //Processor 131 control and data signals
	wire wrProc131West;
	wire fullProc131West;
	wire [31:0] dataOutProc131West;

	//Processor 132 control and data signals
	wire rdProc132North;
	wire emptyProc132North;
	wire [31:0] dataInProc132North;

	 //Processor 132 control and data signals
	wire wrProc132North;
	wire fullProc132North;
	wire [31:0] dataOutProc132North;

	 //Processor 132 control and data signals
	wire rdProc132South;
	wire emptyProc132South;
	wire [31:0] dataInProc132South;
	
	 //Processor 132 control and data signals
	wire wrProc132South;
	wire fullProc132South;
	wire [31:0] dataOutProc132South;

	 //Processor 132 control and data signals
	wire rdProc132East;
	wire emptyProc132East;
	wire [31:0] dataInProc132East;
	
	 //Processor 132 control and data signals
	wire wrProc132East;
	wire fullProc132East;
	wire [31:0] dataOutProc132East;

	 //Processor 132 control and data signals
	wire rdProc132West;
	wire emptyProc132West;
	wire [31:0] dataInProc132West;

	 //Processor 132 control and data signals
	wire wrProc132West;
	wire fullProc132West;
	wire [31:0] dataOutProc132West;

	//Processor 133 control and data signals
	wire rdProc133North;
	wire emptyProc133North;
	wire [31:0] dataInProc133North;

	 //Processor 133 control and data signals
	wire wrProc133North;
	wire fullProc133North;
	wire [31:0] dataOutProc133North;

	 //Processor 133 control and data signals
	wire rdProc133South;
	wire emptyProc133South;
	wire [31:0] dataInProc133South;
	
	 //Processor 133 control and data signals
	wire wrProc133South;
	wire fullProc133South;
	wire [31:0] dataOutProc133South;

	 //Processor 133 control and data signals
	wire rdProc133East;
	wire emptyProc133East;
	wire [31:0] dataInProc133East;
	
	 //Processor 133 control and data signals
	wire wrProc133East;
	wire fullProc133East;
	wire [31:0] dataOutProc133East;

	 //Processor 133 control and data signals
	wire rdProc133West;
	wire emptyProc133West;
	wire [31:0] dataInProc133West;

	 //Processor 133 control and data signals
	wire wrProc133West;
	wire fullProc133West;
	wire [31:0] dataOutProc133West;

	//Processor 134 control and data signals
	wire rdProc134North;
	wire emptyProc134North;
	wire [31:0] dataInProc134North;

	 //Processor 134 control and data signals
	wire wrProc134North;
	wire fullProc134North;
	wire [31:0] dataOutProc134North;

	 //Processor 134 control and data signals
	wire rdProc134South;
	wire emptyProc134South;
	wire [31:0] dataInProc134South;
	
	 //Processor 134 control and data signals
	wire wrProc134South;
	wire fullProc134South;
	wire [31:0] dataOutProc134South;

	 //Processor 134 control and data signals
	wire rdProc134East;
	wire emptyProc134East;
	wire [31:0] dataInProc134East;
	
	 //Processor 134 control and data signals
	wire wrProc134East;
	wire fullProc134East;
	wire [31:0] dataOutProc134East;

	 //Processor 134 control and data signals
	wire rdProc134West;
	wire emptyProc134West;
	wire [31:0] dataInProc134West;

	 //Processor 134 control and data signals
	wire wrProc134West;
	wire fullProc134West;
	wire [31:0] dataOutProc134West;

	//Processor 135 control and data signals
	wire rdProc135North;
	wire emptyProc135North;
	wire [31:0] dataInProc135North;

	 //Processor 135 control and data signals
	wire wrProc135North;
	wire fullProc135North;
	wire [31:0] dataOutProc135North;

	 //Processor 135 control and data signals
	wire rdProc135South;
	wire emptyProc135South;
	wire [31:0] dataInProc135South;
	
	 //Processor 135 control and data signals
	wire wrProc135South;
	wire fullProc135South;
	wire [31:0] dataOutProc135South;

	 //Processor 135 control and data signals
	wire rdProc135East;
	wire emptyProc135East;
	wire [31:0] dataInProc135East;
	
	 //Processor 135 control and data signals
	wire wrProc135East;
	wire fullProc135East;
	wire [31:0] dataOutProc135East;

	 //Processor 135 control and data signals
	wire rdProc135West;
	wire emptyProc135West;
	wire [31:0] dataInProc135West;

	 //Processor 135 control and data signals
	wire wrProc135West;
	wire fullProc135West;
	wire [31:0] dataOutProc135West;

	//Processor 136 control and data signals
	wire rdProc136North;
	wire emptyProc136North;
	wire [31:0] dataInProc136North;

	 //Processor 136 control and data signals
	wire wrProc136North;
	wire fullProc136North;
	wire [31:0] dataOutProc136North;

	 //Processor 136 control and data signals
	wire rdProc136South;
	wire emptyProc136South;
	wire [31:0] dataInProc136South;
	
	 //Processor 136 control and data signals
	wire wrProc136South;
	wire fullProc136South;
	wire [31:0] dataOutProc136South;

	 //Processor 136 control and data signals
	wire rdProc136East;
	wire emptyProc136East;
	wire [31:0] dataInProc136East;
	
	 //Processor 136 control and data signals
	wire wrProc136East;
	wire fullProc136East;
	wire [31:0] dataOutProc136East;

	 //Processor 136 control and data signals
	wire rdProc136West;
	wire emptyProc136West;
	wire [31:0] dataInProc136West;

	 //Processor 136 control and data signals
	wire wrProc136West;
	wire fullProc136West;
	wire [31:0] dataOutProc136West;

	//Processor 137 control and data signals
	wire rdProc137North;
	wire emptyProc137North;
	wire [31:0] dataInProc137North;

	 //Processor 137 control and data signals
	wire wrProc137North;
	wire fullProc137North;
	wire [31:0] dataOutProc137North;

	 //Processor 137 control and data signals
	wire rdProc137South;
	wire emptyProc137South;
	wire [31:0] dataInProc137South;
	
	 //Processor 137 control and data signals
	wire wrProc137South;
	wire fullProc137South;
	wire [31:0] dataOutProc137South;

	 //Processor 137 control and data signals
	wire rdProc137East;
	wire emptyProc137East;
	wire [31:0] dataInProc137East;
	
	 //Processor 137 control and data signals
	wire wrProc137East;
	wire fullProc137East;
	wire [31:0] dataOutProc137East;

	 //Processor 137 control and data signals
	wire rdProc137West;
	wire emptyProc137West;
	wire [31:0] dataInProc137West;

	 //Processor 137 control and data signals
	wire wrProc137West;
	wire fullProc137West;
	wire [31:0] dataOutProc137West;

	//Processor 138 control and data signals
	wire rdProc138North;
	wire emptyProc138North;
	wire [31:0] dataInProc138North;

	 //Processor 138 control and data signals
	wire wrProc138North;
	wire fullProc138North;
	wire [31:0] dataOutProc138North;

	 //Processor 138 control and data signals
	wire rdProc138South;
	wire emptyProc138South;
	wire [31:0] dataInProc138South;
	
	 //Processor 138 control and data signals
	wire wrProc138South;
	wire fullProc138South;
	wire [31:0] dataOutProc138South;

	 //Processor 138 control and data signals
	wire rdProc138East;
	wire emptyProc138East;
	wire [31:0] dataInProc138East;
	
	 //Processor 138 control and data signals
	wire wrProc138East;
	wire fullProc138East;
	wire [31:0] dataOutProc138East;

	 //Processor 138 control and data signals
	wire rdProc138West;
	wire emptyProc138West;
	wire [31:0] dataInProc138West;

	 //Processor 138 control and data signals
	wire wrProc138West;
	wire fullProc138West;
	wire [31:0] dataOutProc138West;

	//Processor 139 control and data signals
	wire rdProc139North;
	wire emptyProc139North;
	wire [31:0] dataInProc139North;

	 //Processor 139 control and data signals
	wire wrProc139North;
	wire fullProc139North;
	wire [31:0] dataOutProc139North;

	 //Processor 139 control and data signals
	wire rdProc139South;
	wire emptyProc139South;
	wire [31:0] dataInProc139South;
	
	 //Processor 139 control and data signals
	wire wrProc139South;
	wire fullProc139South;
	wire [31:0] dataOutProc139South;

	 //Processor 139 control and data signals
	wire rdProc139East;
	wire emptyProc139East;
	wire [31:0] dataInProc139East;
	
	 //Processor 139 control and data signals
	wire wrProc139East;
	wire fullProc139East;
	wire [31:0] dataOutProc139East;

	 //Processor 139 control and data signals
	wire rdProc139West;
	wire emptyProc139West;
	wire [31:0] dataInProc139West;

	 //Processor 139 control and data signals
	wire wrProc139West;
	wire fullProc139West;
	wire [31:0] dataOutProc139West;

	//Processor 140 control and data signals
	wire rdProc140North;
	wire emptyProc140North;
	wire [31:0] dataInProc140North;

	 //Processor 140 control and data signals
	wire wrProc140North;
	wire fullProc140North;
	wire [31:0] dataOutProc140North;

	 //Processor 140 control and data signals
	wire rdProc140South;
	wire emptyProc140South;
	wire [31:0] dataInProc140South;
	
	 //Processor 140 control and data signals
	wire wrProc140South;
	wire fullProc140South;
	wire [31:0] dataOutProc140South;

	 //Processor 140 control and data signals
	wire rdProc140East;
	wire emptyProc140East;
	wire [31:0] dataInProc140East;
	
	 //Processor 140 control and data signals
	wire wrProc140East;
	wire fullProc140East;
	wire [31:0] dataOutProc140East;

	 //Processor 140 control and data signals
	wire rdProc140West;
	wire emptyProc140West;
	wire [31:0] dataInProc140West;

	 //Processor 140 control and data signals
	wire wrProc140West;
	wire fullProc140West;
	wire [31:0] dataOutProc140West;

	//Processor 141 control and data signals
	wire rdProc141North;
	wire emptyProc141North;
	wire [31:0] dataInProc141North;

	 //Processor 141 control and data signals
	wire wrProc141North;
	wire fullProc141North;
	wire [31:0] dataOutProc141North;

	 //Processor 141 control and data signals
	wire rdProc141South;
	wire emptyProc141South;
	wire [31:0] dataInProc141South;
	
	 //Processor 141 control and data signals
	wire wrProc141South;
	wire fullProc141South;
	wire [31:0] dataOutProc141South;

	 //Processor 141 control and data signals
	wire rdProc141East;
	wire emptyProc141East;
	wire [31:0] dataInProc141East;
	
	 //Processor 141 control and data signals
	wire wrProc141East;
	wire fullProc141East;
	wire [31:0] dataOutProc141East;

	 //Processor 141 control and data signals
	wire rdProc141West;
	wire emptyProc141West;
	wire [31:0] dataInProc141West;

	 //Processor 141 control and data signals
	wire wrProc141West;
	wire fullProc141West;
	wire [31:0] dataOutProc141West;

	//Processor 142 control and data signals
	wire wrProc142North;
	wire fullProc142North;
	wire [31:0] dataOutProc142North;

	//Processor 142 control and data signals
        wire rdProc142North;
        wire emptyProc142North;
        wire [31:0] dataInProc142North;

	//Processor 142 control and data signals
	wire rdProc142South;
	wire emptyProc142South;
	wire [31:0] dataInProc142South;
		
	 //Processor 142 control and data signals
	wire wrProc142South;
	wire fullProc142South;
	wire [31:0] dataOutProc142South;

	 //Processor 142 control and data signals
	wire wrProc142West;
	wire fullProc142West;
	wire [31:0] dataOutProc142West;
	
	 //Processor 142 control and data signals
	wire rdProc142West;
	wire emptyProc142West;
	wire [31:0] dataInProc142West;

	 //Processor143 control and data signals
	wire wrProc143North;
	wire fullProc143North;
	wire [31:0] dataOutProc143North;
	
	 //Processor 143 control and data signals
	wire rdProc143North;
	wire emptyProc143North;
	wire [31:0] dataInProc143North;

	 //Processor 143 control and data signals
	wire rdProc143East;
	wire emptyProc143East;
	wire [31:0] dataInProc143East;

	 //Processor 143 control and data signals
	wire wrProc143East;
	wire fullProc143East;
	wire [31:0] dataOutProc143East;

	//Processor 144 control and data signals
	wire wrProc144North;
	wire fullProc144North;
	wire [31:0] dataOutProc144North;
		
	 //Processor 144 control and data signals
	wire rdProc144North;
	wire emptyProc144North;
	wire [31:0] dataInProc144North;

	 //Processor 144 control and data signals
	wire rdProc144East;
	wire emptyProc144East;
	wire [31:0] dataInProc144East;
	
	 //Processor 144 control and data signals
	wire wrProc144East;
	wire fullProc144East;
	wire [31:0] dataOutProc144East;

	 //Processor 144 control and data signals
	wire rdProc144West;
	wire emptyProc144West;
	wire [31:0] dataInProc144West;

	 //Processor 144 control and data signals
	wire wrProc144West;
	wire fullProc144West;
	wire [31:0] dataOutProc144West;

	//Processor 145 control and data signals
	wire wrProc145North;
	wire fullProc145North;
	wire [31:0] dataOutProc145North;
		
	 //Processor 145 control and data signals
	wire rdProc145North;
	wire emptyProc145North;
	wire [31:0] dataInProc145North;

	 //Processor 145 control and data signals
	wire rdProc145East;
	wire emptyProc145East;
	wire [31:0] dataInProc145East;
	
	 //Processor 145 control and data signals
	wire wrProc145East;
	wire fullProc145East;
	wire [31:0] dataOutProc145East;

	 //Processor 145 control and data signals
	wire rdProc145West;
	wire emptyProc145West;
	wire [31:0] dataInProc145West;

	 //Processor 145 control and data signals
	wire wrProc145West;
	wire fullProc145West;
	wire [31:0] dataOutProc145West;

	//Processor 146 control and data signals
	wire wrProc146North;
	wire fullProc146North;
	wire [31:0] dataOutProc146North;
		
	 //Processor 146 control and data signals
	wire rdProc146North;
	wire emptyProc146North;
	wire [31:0] dataInProc146North;

	 //Processor 146 control and data signals
	wire rdProc146East;
	wire emptyProc146East;
	wire [31:0] dataInProc146East;
	
	 //Processor 146 control and data signals
	wire wrProc146East;
	wire fullProc146East;
	wire [31:0] dataOutProc146East;

	 //Processor 146 control and data signals
	wire rdProc146West;
	wire emptyProc146West;
	wire [31:0] dataInProc146West;

	 //Processor 146 control and data signals
	wire wrProc146West;
	wire fullProc146West;
	wire [31:0] dataOutProc146West;

	//Processor 147 control and data signals
	wire wrProc147North;
	wire fullProc147North;
	wire [31:0] dataOutProc147North;
		
	 //Processor 147 control and data signals
	wire rdProc147North;
	wire emptyProc147North;
	wire [31:0] dataInProc147North;

	 //Processor 147 control and data signals
	wire rdProc147East;
	wire emptyProc147East;
	wire [31:0] dataInProc147East;
	
	 //Processor 147 control and data signals
	wire wrProc147East;
	wire fullProc147East;
	wire [31:0] dataOutProc147East;

	 //Processor 147 control and data signals
	wire rdProc147West;
	wire emptyProc147West;
	wire [31:0] dataInProc147West;

	 //Processor 147 control and data signals
	wire wrProc147West;
	wire fullProc147West;
	wire [31:0] dataOutProc147West;

	//Processor 148 control and data signals
	wire wrProc148North;
	wire fullProc148North;
	wire [31:0] dataOutProc148North;
		
	 //Processor 148 control and data signals
	wire rdProc148North;
	wire emptyProc148North;
	wire [31:0] dataInProc148North;

	 //Processor 148 control and data signals
	wire rdProc148East;
	wire emptyProc148East;
	wire [31:0] dataInProc148East;
	
	 //Processor 148 control and data signals
	wire wrProc148East;
	wire fullProc148East;
	wire [31:0] dataOutProc148East;

	 //Processor 148 control and data signals
	wire rdProc148West;
	wire emptyProc148West;
	wire [31:0] dataInProc148West;

	 //Processor 148 control and data signals
	wire wrProc148West;
	wire fullProc148West;
	wire [31:0] dataOutProc148West;

	//Processor 149 control and data signals
	wire wrProc149North;
	wire fullProc149North;
	wire [31:0] dataOutProc149North;
		
	 //Processor 149 control and data signals
	wire rdProc149North;
	wire emptyProc149North;
	wire [31:0] dataInProc149North;

	 //Processor 149 control and data signals
	wire rdProc149East;
	wire emptyProc149East;
	wire [31:0] dataInProc149East;
	
	 //Processor 149 control and data signals
	wire wrProc149East;
	wire fullProc149East;
	wire [31:0] dataOutProc149East;

	 //Processor 149 control and data signals
	wire rdProc149West;
	wire emptyProc149West;
	wire [31:0] dataInProc149West;

	 //Processor 149 control and data signals
	wire wrProc149West;
	wire fullProc149West;
	wire [31:0] dataOutProc149West;

	//Processor 150 control and data signals
	wire wrProc150North;
	wire fullProc150North;
	wire [31:0] dataOutProc150North;
		
	 //Processor 150 control and data signals
	wire rdProc150North;
	wire emptyProc150North;
	wire [31:0] dataInProc150North;

	 //Processor 150 control and data signals
	wire rdProc150East;
	wire emptyProc150East;
	wire [31:0] dataInProc150East;
	
	 //Processor 150 control and data signals
	wire wrProc150East;
	wire fullProc150East;
	wire [31:0] dataOutProc150East;

	 //Processor 150 control and data signals
	wire rdProc150West;
	wire emptyProc150West;
	wire [31:0] dataInProc150West;

	 //Processor 150 control and data signals
	wire wrProc150West;
	wire fullProc150West;
	wire [31:0] dataOutProc150West;

	//Processor 151 control and data signals
	wire wrProc151North;
	wire fullProc151North;
	wire [31:0] dataOutProc151North;
		
	 //Processor 151 control and data signals
	wire rdProc151North;
	wire emptyProc151North;
	wire [31:0] dataInProc151North;

	 //Processor 151 control and data signals
	wire rdProc151East;
	wire emptyProc151East;
	wire [31:0] dataInProc151East;
	
	 //Processor 151 control and data signals
	wire wrProc151East;
	wire fullProc151East;
	wire [31:0] dataOutProc151East;

	 //Processor 151 control and data signals
	wire rdProc151West;
	wire emptyProc151West;
	wire [31:0] dataInProc151West;

	 //Processor 151 control and data signals
	wire wrProc151West;
	wire fullProc151West;
	wire [31:0] dataOutProc151West;

	//Processor 152 control and data signals
	wire wrProc152North;
	wire fullProc152North;
	wire [31:0] dataOutProc152North;
		
	 //Processor 152 control and data signals
	wire rdProc152North;
	wire emptyProc152North;
	wire [31:0] dataInProc152North;

	 //Processor 152 control and data signals
	wire rdProc152East;
	wire emptyProc152East;
	wire [31:0] dataInProc152East;
	
	 //Processor 152 control and data signals
	wire wrProc152East;
	wire fullProc152East;
	wire [31:0] dataOutProc152East;

	 //Processor 152 control and data signals
	wire rdProc152West;
	wire emptyProc152West;
	wire [31:0] dataInProc152West;

	 //Processor 152 control and data signals
	wire wrProc152West;
	wire fullProc152West;
	wire [31:0] dataOutProc152West;

	//Processor 153 control and data signals
	wire wrProc153North;
	wire fullProc153North;
	wire [31:0] dataOutProc153North;
		
	 //Processor 153 control and data signals
	wire rdProc153North;
	wire emptyProc153North;
	wire [31:0] dataInProc153North;

	 //Processor 153 control and data signals
	wire rdProc153East;
	wire emptyProc153East;
	wire [31:0] dataInProc153East;
	
	 //Processor 153 control and data signals
	wire wrProc153East;
	wire fullProc153East;
	wire [31:0] dataOutProc153East;

	 //Processor 153 control and data signals
	wire rdProc153West;
	wire emptyProc153West;
	wire [31:0] dataInProc153West;

	 //Processor 153 control and data signals
	wire wrProc153West;
	wire fullProc153West;
	wire [31:0] dataOutProc153West;

	//Processor 154 control and data signals
	wire wrProc154North;
	wire fullProc154North;
	wire [31:0] dataOutProc154North;
		
	 //Processor 154 control and data signals
	wire rdProc154North;
	wire emptyProc154North;
	wire [31:0] dataInProc154North;

	 //Processor 154 control and data signals
	wire rdProc154East;
	wire emptyProc154East;
	wire [31:0] dataInProc154East;
	
	 //Processor 154 control and data signals
	wire wrProc154East;
	wire fullProc154East;
	wire [31:0] dataOutProc154East;

	 //Processor 154 control and data signals
	wire rdProc154West;
	wire emptyProc154West;
	wire [31:0] dataInProc154West;

	 //Processor 154 control and data signals
	wire wrProc154West;
	wire fullProc154West;
	wire [31:0] dataOutProc154West;

	//Processor 155 control and data signals
	wire rdProc155North;
	wire emptyProc155North;
	wire [31:0] dataInProc155North;

	 //Processor 155 control and data signals
	wire wrProc155North;
	wire fullProc155North;
	wire [31:0] dataOutProc155North;

	 //Processor 155 control and data signals
	wire wrProc155West;
	wire fullProc155West;
	wire [31:0] dataOutProc155West;
	
	 //Processor 155 control and data signals
	wire rdProc155West;
	wire emptyProc155West;
	wire [31:0] dataInProc155West;

 
//PROCESSOR 0
system proc0(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe0),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe0),
	.rdSouth(rdProc0South),
	.emptySouth(emptyProc0South),
	.dataInSouth(dataInProc0South),
	.wrSouth(wrProc0South),
	.fullSouth(fullProc0South),
	.dataOutSouth(dataOutProc0South),
	.rdEast(rdProc0East),
	.emptyEast(emptyProc0East),
	.dataInEast(dataInProc0East),
	.wrEast(wrProc0East),
	.fullEast(fullProc0East),
	.dataOutEast(dataOutProc0East),

	.reg_file_b_readdataout(reg_file_b_readdataout));
 
//PROCESSOR 1
system proc1(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe1),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe1),	
	.rdSouth(rdProc1South),
	.emptySouth(emptyProc1South),
	.dataInSouth(dataInProc1South),
	.wrSouth(wrProc1South),
	.fullSouth(fullProc1South),
	.dataOutSouth(dataOutProc1South),
	.rdEast(rdProc1East),
	.emptyEast(emptyProc1East),
	.dataInEast(dataInProc1East),
	.wrEast(wrProc1East),
	.fullEast(fullProc1East),
	.dataOutEast(dataOutProc1East),
	.rdWest(rdProc1West),
	.emptyWest(emptyProc1West),
	.dataInWest(dataInProc1West),
	.wrWest(wrProc1West),
	.fullWest(fullProc1West),
	.dataOutWest(dataOutProc1West));
 
//PROCESSOR 2
system proc2(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe2),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe2),	
	.rdSouth(rdProc2South),
	.emptySouth(emptyProc2South),
	.dataInSouth(dataInProc2South),
	.wrSouth(wrProc2South),
	.fullSouth(fullProc2South),
	.dataOutSouth(dataOutProc2South),
	.rdEast(rdProc2East),
	.emptyEast(emptyProc2East),
	.dataInEast(dataInProc2East),
	.wrEast(wrProc2East),
	.fullEast(fullProc2East),
	.dataOutEast(dataOutProc2East),
	.rdWest(rdProc2West),
	.emptyWest(emptyProc2West),
	.dataInWest(dataInProc2West),
	.wrWest(wrProc2West),
	.fullWest(fullProc2West),
	.dataOutWest(dataOutProc2West));
 
//PROCESSOR 3
system proc3(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe3),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe3),	
	.rdSouth(rdProc3South),
	.emptySouth(emptyProc3South),
	.dataInSouth(dataInProc3South),
	.wrSouth(wrProc3South),
	.fullSouth(fullProc3South),
	.dataOutSouth(dataOutProc3South),
	.rdEast(rdProc3East),
	.emptyEast(emptyProc3East),
	.dataInEast(dataInProc3East),
	.wrEast(wrProc3East),
	.fullEast(fullProc3East),
	.dataOutEast(dataOutProc3East),
	.rdWest(rdProc3West),
	.emptyWest(emptyProc3West),
	.dataInWest(dataInProc3West),
	.wrWest(wrProc3West),
	.fullWest(fullProc3West),
	.dataOutWest(dataOutProc3West));
 
//PROCESSOR 4
system proc4(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe4),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe4),	
	.rdSouth(rdProc4South),
	.emptySouth(emptyProc4South),
	.dataInSouth(dataInProc4South),
	.wrSouth(wrProc4South),
	.fullSouth(fullProc4South),
	.dataOutSouth(dataOutProc4South),
	.rdEast(rdProc4East),
	.emptyEast(emptyProc4East),
	.dataInEast(dataInProc4East),
	.wrEast(wrProc4East),
	.fullEast(fullProc4East),
	.dataOutEast(dataOutProc4East),
	.rdWest(rdProc4West),
	.emptyWest(emptyProc4West),
	.dataInWest(dataInProc4West),
	.wrWest(wrProc4West),
	.fullWest(fullProc4West),
	.dataOutWest(dataOutProc4West));
 
//PROCESSOR 5
system proc5(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe5),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe5),	
	.rdSouth(rdProc5South),
	.emptySouth(emptyProc5South),
	.dataInSouth(dataInProc5South),
	.wrSouth(wrProc5South),
	.fullSouth(fullProc5South),
	.dataOutSouth(dataOutProc5South),
	.rdEast(rdProc5East),
	.emptyEast(emptyProc5East),
	.dataInEast(dataInProc5East),
	.wrEast(wrProc5East),
	.fullEast(fullProc5East),
	.dataOutEast(dataOutProc5East),
	.rdWest(rdProc5West),
	.emptyWest(emptyProc5West),
	.dataInWest(dataInProc5West),
	.wrWest(wrProc5West),
	.fullWest(fullProc5West),
	.dataOutWest(dataOutProc5West));
 
//PROCESSOR 6
system proc6(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe6),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe6),	
	.rdSouth(rdProc6South),
	.emptySouth(emptyProc6South),
	.dataInSouth(dataInProc6South),
	.wrSouth(wrProc6South),
	.fullSouth(fullProc6South),
	.dataOutSouth(dataOutProc6South),
	.rdEast(rdProc6East),
	.emptyEast(emptyProc6East),
	.dataInEast(dataInProc6East),
	.wrEast(wrProc6East),
	.fullEast(fullProc6East),
	.dataOutEast(dataOutProc6East),
	.rdWest(rdProc6West),
	.emptyWest(emptyProc6West),
	.dataInWest(dataInProc6West),
	.wrWest(wrProc6West),
	.fullWest(fullProc6West),
	.dataOutWest(dataOutProc6West));
 
//PROCESSOR 7
system proc7(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe7),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe7),	
	.rdSouth(rdProc7South),
	.emptySouth(emptyProc7South),
	.dataInSouth(dataInProc7South),
	.wrSouth(wrProc7South),
	.fullSouth(fullProc7South),
	.dataOutSouth(dataOutProc7South),
	.rdEast(rdProc7East),
	.emptyEast(emptyProc7East),
	.dataInEast(dataInProc7East),
	.wrEast(wrProc7East),
	.fullEast(fullProc7East),
	.dataOutEast(dataOutProc7East),
	.rdWest(rdProc7West),
	.emptyWest(emptyProc7West),
	.dataInWest(dataInProc7West),
	.wrWest(wrProc7West),
	.fullWest(fullProc7West),
	.dataOutWest(dataOutProc7West));
 
//PROCESSOR 8
system proc8(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe8),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe8),	
	.rdSouth(rdProc8South),
	.emptySouth(emptyProc8South),
	.dataInSouth(dataInProc8South),
	.wrSouth(wrProc8South),
	.fullSouth(fullProc8South),
	.dataOutSouth(dataOutProc8South),
	.rdEast(rdProc8East),
	.emptyEast(emptyProc8East),
	.dataInEast(dataInProc8East),
	.wrEast(wrProc8East),
	.fullEast(fullProc8East),
	.dataOutEast(dataOutProc8East),
	.rdWest(rdProc8West),
	.emptyWest(emptyProc8West),
	.dataInWest(dataInProc8West),
	.wrWest(wrProc8West),
	.fullWest(fullProc8West),
	.dataOutWest(dataOutProc8West));
 
//PROCESSOR 9
system proc9(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe9),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe9),	
	.rdSouth(rdProc9South),
	.emptySouth(emptyProc9South),
	.dataInSouth(dataInProc9South),
	.wrSouth(wrProc9South),
	.fullSouth(fullProc9South),
	.dataOutSouth(dataOutProc9South),
	.rdEast(rdProc9East),
	.emptyEast(emptyProc9East),
	.dataInEast(dataInProc9East),
	.wrEast(wrProc9East),
	.fullEast(fullProc9East),
	.dataOutEast(dataOutProc9East),
	.rdWest(rdProc9West),
	.emptyWest(emptyProc9West),
	.dataInWest(dataInProc9West),
	.wrWest(wrProc9West),
	.fullWest(fullProc9West),
	.dataOutWest(dataOutProc9West));
 
//PROCESSOR 10
system proc10(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe10),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe10),	
	.rdSouth(rdProc10South),
	.emptySouth(emptyProc10South),
	.dataInSouth(dataInProc10South),
	.wrSouth(wrProc10South),
	.fullSouth(fullProc10South),
	.dataOutSouth(dataOutProc10South),
	.rdEast(rdProc10East),
	.emptyEast(emptyProc10East),
	.dataInEast(dataInProc10East),
	.wrEast(wrProc10East),
	.fullEast(fullProc10East),
	.dataOutEast(dataOutProc10East),
	.rdWest(rdProc10West),
	.emptyWest(emptyProc10West),
	.dataInWest(dataInProc10West),
	.wrWest(wrProc10West),
	.fullWest(fullProc10West),
	.dataOutWest(dataOutProc10West));
 
//PROCESSOR 11
system proc11(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe11),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe11),	
	.rdSouth(rdProc11South),
	.emptySouth(emptyProc11South),
	.dataInSouth(dataInProc11South),
	.wrSouth(wrProc11South),
	.fullSouth(fullProc11South),
	.dataOutSouth(dataOutProc11South),
	.rdEast(rdProc11East),
	.emptyEast(emptyProc11East),
	.dataInEast(dataInProc11East),
	.wrEast(wrProc11East),
	.fullEast(fullProc11East),
	.dataOutEast(dataOutProc11East),
	.rdWest(rdProc11West),
	.emptyWest(emptyProc11West),
	.dataInWest(dataInProc11West),
	.wrWest(wrProc11West),
	.fullWest(fullProc11West),
	.dataOutWest(dataOutProc11West));
 
//PROCESSOR 12
system proc12(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe12),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe12),	
	.rdSouth(rdProc12South),
	.emptySouth(emptyProc12South),
	.dataInSouth(dataInProc12South),
	.wrSouth(wrProc12South),
	.fullSouth(fullProc12South),
	.dataOutSouth(dataOutProc12South),
	.rdWest(rdProc12West),
	.emptyWest(emptyProc12West),
	.dataInWest(dataInProc12West),
	.wrWest(wrProc12West),
	.fullWest(fullProc12West),
	.dataOutWest(dataOutProc12West));
 
//PROCESSOR 13
system proc13(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe13),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe13),
	.wrNorth(wrProc13North),
	.fullNorth(fullProc13North),
	.dataOutNorth(dataOutProc13North),
	.rdNorth(rdProc13North),
	.emptyNorth(emptyProc13North),
	.dataInNorth(dataInProc13North),
	.rdSouth(rdProc13South),
	.emptySouth(emptyProc13South),
	.dataInSouth(dataInProc13South),
	.wrSouth(wrProc13South),
	.fullSouth(fullProc13South),
	.dataOutSouth(dataOutProc13South),
	.rdEast(rdProc13East),
	.emptyEast(emptyProc13East),
	.dataInEast(dataInProc13East),
	.wrEast(wrProc13East),
	.fullEast(fullProc13East),
	.dataOutEast(dataOutProc13East));
 
//PROCESSOR 14
system proc14(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe14),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe14),
	.rdNorth(rdProc14North),
	.emptyNorth(emptyProc14North),
	.dataInNorth(dataInProc14North),
	.wrNorth(wrProc14North),
	.fullNorth(fullProc14North),
	.dataOutNorth(dataOutProc14North),
	.rdSouth(rdProc14South),
	.emptySouth(emptyProc14South),
	.dataInSouth(dataInProc14South),
	.wrSouth(wrProc14South),
	.fullSouth(fullProc14South),
	.dataOutSouth(dataOutProc14South),
	.rdEast(rdProc14East),
	.emptyEast(emptyProc14East),
	.dataInEast(dataInProc14East),
	.wrEast(wrProc14East),
	.fullEast(fullProc14East),
	.dataOutEast(dataOutProc14East),
	.rdWest(rdProc14West),
	.emptyWest(emptyProc14West),
	.dataInWest(dataInProc14West),
	.wrWest(wrProc14West),
	.fullWest(fullProc14West),
	.dataOutWest(dataOutProc14West));
 
//PROCESSOR 15
system proc15(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe15),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe15),
	.rdNorth(rdProc15North),
	.emptyNorth(emptyProc15North),
	.dataInNorth(dataInProc15North),
	.wrNorth(wrProc15North),
	.fullNorth(fullProc15North),
	.dataOutNorth(dataOutProc15North),
	.rdSouth(rdProc15South),
	.emptySouth(emptyProc15South),
	.dataInSouth(dataInProc15South),
	.wrSouth(wrProc15South),
	.fullSouth(fullProc15South),
	.dataOutSouth(dataOutProc15South),
	.rdEast(rdProc15East),
	.emptyEast(emptyProc15East),
	.dataInEast(dataInProc15East),
	.wrEast(wrProc15East),
	.fullEast(fullProc15East),
	.dataOutEast(dataOutProc15East),
	.rdWest(rdProc15West),
	.emptyWest(emptyProc15West),
	.dataInWest(dataInProc15West),
	.wrWest(wrProc15West),
	.fullWest(fullProc15West),
	.dataOutWest(dataOutProc15West));
 
//PROCESSOR 16
system proc16(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe16),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe16),
	.rdNorth(rdProc16North),
	.emptyNorth(emptyProc16North),
	.dataInNorth(dataInProc16North),
	.wrNorth(wrProc16North),
	.fullNorth(fullProc16North),
	.dataOutNorth(dataOutProc16North),
	.rdSouth(rdProc16South),
	.emptySouth(emptyProc16South),
	.dataInSouth(dataInProc16South),
	.wrSouth(wrProc16South),
	.fullSouth(fullProc16South),
	.dataOutSouth(dataOutProc16South),
	.rdEast(rdProc16East),
	.emptyEast(emptyProc16East),
	.dataInEast(dataInProc16East),
	.wrEast(wrProc16East),
	.fullEast(fullProc16East),
	.dataOutEast(dataOutProc16East),
	.rdWest(rdProc16West),
	.emptyWest(emptyProc16West),
	.dataInWest(dataInProc16West),
	.wrWest(wrProc16West),
	.fullWest(fullProc16West),
	.dataOutWest(dataOutProc16West));
 
//PROCESSOR 17
system proc17(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe17),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe17),
	.rdNorth(rdProc17North),
	.emptyNorth(emptyProc17North),
	.dataInNorth(dataInProc17North),
	.wrNorth(wrProc17North),
	.fullNorth(fullProc17North),
	.dataOutNorth(dataOutProc17North),
	.rdSouth(rdProc17South),
	.emptySouth(emptyProc17South),
	.dataInSouth(dataInProc17South),
	.wrSouth(wrProc17South),
	.fullSouth(fullProc17South),
	.dataOutSouth(dataOutProc17South),
	.rdEast(rdProc17East),
	.emptyEast(emptyProc17East),
	.dataInEast(dataInProc17East),
	.wrEast(wrProc17East),
	.fullEast(fullProc17East),
	.dataOutEast(dataOutProc17East),
	.rdWest(rdProc17West),
	.emptyWest(emptyProc17West),
	.dataInWest(dataInProc17West),
	.wrWest(wrProc17West),
	.fullWest(fullProc17West),
	.dataOutWest(dataOutProc17West));
 
//PROCESSOR 18
system proc18(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe18),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe18),
	.rdNorth(rdProc18North),
	.emptyNorth(emptyProc18North),
	.dataInNorth(dataInProc18North),
	.wrNorth(wrProc18North),
	.fullNorth(fullProc18North),
	.dataOutNorth(dataOutProc18North),
	.rdSouth(rdProc18South),
	.emptySouth(emptyProc18South),
	.dataInSouth(dataInProc18South),
	.wrSouth(wrProc18South),
	.fullSouth(fullProc18South),
	.dataOutSouth(dataOutProc18South),
	.rdEast(rdProc18East),
	.emptyEast(emptyProc18East),
	.dataInEast(dataInProc18East),
	.wrEast(wrProc18East),
	.fullEast(fullProc18East),
	.dataOutEast(dataOutProc18East),
	.rdWest(rdProc18West),
	.emptyWest(emptyProc18West),
	.dataInWest(dataInProc18West),
	.wrWest(wrProc18West),
	.fullWest(fullProc18West),
	.dataOutWest(dataOutProc18West));
 
//PROCESSOR 19
system proc19(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe19),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe19),
	.rdNorth(rdProc19North),
	.emptyNorth(emptyProc19North),
	.dataInNorth(dataInProc19North),
	.wrNorth(wrProc19North),
	.fullNorth(fullProc19North),
	.dataOutNorth(dataOutProc19North),
	.rdSouth(rdProc19South),
	.emptySouth(emptyProc19South),
	.dataInSouth(dataInProc19South),
	.wrSouth(wrProc19South),
	.fullSouth(fullProc19South),
	.dataOutSouth(dataOutProc19South),
	.rdEast(rdProc19East),
	.emptyEast(emptyProc19East),
	.dataInEast(dataInProc19East),
	.wrEast(wrProc19East),
	.fullEast(fullProc19East),
	.dataOutEast(dataOutProc19East),
	.rdWest(rdProc19West),
	.emptyWest(emptyProc19West),
	.dataInWest(dataInProc19West),
	.wrWest(wrProc19West),
	.fullWest(fullProc19West),
	.dataOutWest(dataOutProc19West));
 
//PROCESSOR 20
system proc20(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe20),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe20),
	.rdNorth(rdProc20North),
	.emptyNorth(emptyProc20North),
	.dataInNorth(dataInProc20North),
	.wrNorth(wrProc20North),
	.fullNorth(fullProc20North),
	.dataOutNorth(dataOutProc20North),
	.rdSouth(rdProc20South),
	.emptySouth(emptyProc20South),
	.dataInSouth(dataInProc20South),
	.wrSouth(wrProc20South),
	.fullSouth(fullProc20South),
	.dataOutSouth(dataOutProc20South),
	.rdEast(rdProc20East),
	.emptyEast(emptyProc20East),
	.dataInEast(dataInProc20East),
	.wrEast(wrProc20East),
	.fullEast(fullProc20East),
	.dataOutEast(dataOutProc20East),
	.rdWest(rdProc20West),
	.emptyWest(emptyProc20West),
	.dataInWest(dataInProc20West),
	.wrWest(wrProc20West),
	.fullWest(fullProc20West),
	.dataOutWest(dataOutProc20West));
 
//PROCESSOR 21
system proc21(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe21),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe21),
	.rdNorth(rdProc21North),
	.emptyNorth(emptyProc21North),
	.dataInNorth(dataInProc21North),
	.wrNorth(wrProc21North),
	.fullNorth(fullProc21North),
	.dataOutNorth(dataOutProc21North),
	.rdSouth(rdProc21South),
	.emptySouth(emptyProc21South),
	.dataInSouth(dataInProc21South),
	.wrSouth(wrProc21South),
	.fullSouth(fullProc21South),
	.dataOutSouth(dataOutProc21South),
	.rdEast(rdProc21East),
	.emptyEast(emptyProc21East),
	.dataInEast(dataInProc21East),
	.wrEast(wrProc21East),
	.fullEast(fullProc21East),
	.dataOutEast(dataOutProc21East),
	.rdWest(rdProc21West),
	.emptyWest(emptyProc21West),
	.dataInWest(dataInProc21West),
	.wrWest(wrProc21West),
	.fullWest(fullProc21West),
	.dataOutWest(dataOutProc21West));
 
//PROCESSOR 22
system proc22(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe22),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe22),
	.rdNorth(rdProc22North),
	.emptyNorth(emptyProc22North),
	.dataInNorth(dataInProc22North),
	.wrNorth(wrProc22North),
	.fullNorth(fullProc22North),
	.dataOutNorth(dataOutProc22North),
	.rdSouth(rdProc22South),
	.emptySouth(emptyProc22South),
	.dataInSouth(dataInProc22South),
	.wrSouth(wrProc22South),
	.fullSouth(fullProc22South),
	.dataOutSouth(dataOutProc22South),
	.rdEast(rdProc22East),
	.emptyEast(emptyProc22East),
	.dataInEast(dataInProc22East),
	.wrEast(wrProc22East),
	.fullEast(fullProc22East),
	.dataOutEast(dataOutProc22East),
	.rdWest(rdProc22West),
	.emptyWest(emptyProc22West),
	.dataInWest(dataInProc22West),
	.wrWest(wrProc22West),
	.fullWest(fullProc22West),
	.dataOutWest(dataOutProc22West));
 
//PROCESSOR 23
system proc23(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe23),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe23),
	.rdNorth(rdProc23North),
	.emptyNorth(emptyProc23North),
	.dataInNorth(dataInProc23North),
	.wrNorth(wrProc23North),
	.fullNorth(fullProc23North),
	.dataOutNorth(dataOutProc23North),
	.rdSouth(rdProc23South),
	.emptySouth(emptyProc23South),
	.dataInSouth(dataInProc23South),
	.wrSouth(wrProc23South),
	.fullSouth(fullProc23South),
	.dataOutSouth(dataOutProc23South),
	.rdEast(rdProc23East),
	.emptyEast(emptyProc23East),
	.dataInEast(dataInProc23East),
	.wrEast(wrProc23East),
	.fullEast(fullProc23East),
	.dataOutEast(dataOutProc23East),
	.rdWest(rdProc23West),
	.emptyWest(emptyProc23West),
	.dataInWest(dataInProc23West),
	.wrWest(wrProc23West),
	.fullWest(fullProc23West),
	.dataOutWest(dataOutProc23West));
 
//PROCESSOR 24
system proc24(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe24),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe24),
	.rdNorth(rdProc24North),
	.emptyNorth(emptyProc24North),
	.dataInNorth(dataInProc24North),
	.wrNorth(wrProc24North),
	.fullNorth(fullProc24North),
	.dataOutNorth(dataOutProc24North),
	.rdSouth(rdProc24South),
	.emptySouth(emptyProc24South),
	.dataInSouth(dataInProc24South),
	.wrSouth(wrProc24South),
	.fullSouth(fullProc24South),
	.dataOutSouth(dataOutProc24South),
	.rdEast(rdProc24East),
	.emptyEast(emptyProc24East),
	.dataInEast(dataInProc24East),
	.wrEast(wrProc24East),
	.fullEast(fullProc24East),
	.dataOutEast(dataOutProc24East),
	.rdWest(rdProc24West),
	.emptyWest(emptyProc24West),
	.dataInWest(dataInProc24West),
	.wrWest(wrProc24West),
	.fullWest(fullProc24West),
	.dataOutWest(dataOutProc24West));
 
//PROCESSOR 25
system proc25(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe25),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe25),
	.rdNorth(rdProc25North),
	.emptyNorth(emptyProc25North),
	.dataInNorth(dataInProc25North),
	.wrNorth(wrProc25North),
	.fullNorth(fullProc25North),
	.dataOutNorth(dataOutProc25North),
	.rdSouth(rdProc25South),
	.emptySouth(emptyProc25South),
	.dataInSouth(dataInProc25South),
	.wrSouth(wrProc25South),
	.fullSouth(fullProc25South),
	.dataOutSouth(dataOutProc25South),
	.rdWest(rdProc25West),
	.emptyWest(emptyProc25West),
	.dataInWest(dataInProc25West),
	.wrWest(wrProc25West),
	.fullWest(fullProc25West),
	.dataOutWest(dataOutProc25West));
 
//PROCESSOR 26
system proc26(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe26),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe26),
	.wrNorth(wrProc26North),
	.fullNorth(fullProc26North),
	.dataOutNorth(dataOutProc26North),
	.rdNorth(rdProc26North),
	.emptyNorth(emptyProc26North),
	.dataInNorth(dataInProc26North),
	.rdSouth(rdProc26South),
	.emptySouth(emptyProc26South),
	.dataInSouth(dataInProc26South),
	.wrSouth(wrProc26South),
	.fullSouth(fullProc26South),
	.dataOutSouth(dataOutProc26South),
	.rdEast(rdProc26East),
	.emptyEast(emptyProc26East),
	.dataInEast(dataInProc26East),
	.wrEast(wrProc26East),
	.fullEast(fullProc26East),
	.dataOutEast(dataOutProc26East));
 
//PROCESSOR 27
system proc27(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe27),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe27),
	.rdNorth(rdProc27North),
	.emptyNorth(emptyProc27North),
	.dataInNorth(dataInProc27North),
	.wrNorth(wrProc27North),
	.fullNorth(fullProc27North),
	.dataOutNorth(dataOutProc27North),
	.rdSouth(rdProc27South),
	.emptySouth(emptyProc27South),
	.dataInSouth(dataInProc27South),
	.wrSouth(wrProc27South),
	.fullSouth(fullProc27South),
	.dataOutSouth(dataOutProc27South),
	.rdEast(rdProc27East),
	.emptyEast(emptyProc27East),
	.dataInEast(dataInProc27East),
	.wrEast(wrProc27East),
	.fullEast(fullProc27East),
	.dataOutEast(dataOutProc27East),
	.rdWest(rdProc27West),
	.emptyWest(emptyProc27West),
	.dataInWest(dataInProc27West),
	.wrWest(wrProc27West),
	.fullWest(fullProc27West),
	.dataOutWest(dataOutProc27West));
 
//PROCESSOR 28
system proc28(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe28),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe28),
	.rdNorth(rdProc28North),
	.emptyNorth(emptyProc28North),
	.dataInNorth(dataInProc28North),
	.wrNorth(wrProc28North),
	.fullNorth(fullProc28North),
	.dataOutNorth(dataOutProc28North),
	.rdSouth(rdProc28South),
	.emptySouth(emptyProc28South),
	.dataInSouth(dataInProc28South),
	.wrSouth(wrProc28South),
	.fullSouth(fullProc28South),
	.dataOutSouth(dataOutProc28South),
	.rdEast(rdProc28East),
	.emptyEast(emptyProc28East),
	.dataInEast(dataInProc28East),
	.wrEast(wrProc28East),
	.fullEast(fullProc28East),
	.dataOutEast(dataOutProc28East),
	.rdWest(rdProc28West),
	.emptyWest(emptyProc28West),
	.dataInWest(dataInProc28West),
	.wrWest(wrProc28West),
	.fullWest(fullProc28West),
	.dataOutWest(dataOutProc28West));
 
//PROCESSOR 29
system proc29(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe29),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe29),
	.rdNorth(rdProc29North),
	.emptyNorth(emptyProc29North),
	.dataInNorth(dataInProc29North),
	.wrNorth(wrProc29North),
	.fullNorth(fullProc29North),
	.dataOutNorth(dataOutProc29North),
	.rdSouth(rdProc29South),
	.emptySouth(emptyProc29South),
	.dataInSouth(dataInProc29South),
	.wrSouth(wrProc29South),
	.fullSouth(fullProc29South),
	.dataOutSouth(dataOutProc29South),
	.rdEast(rdProc29East),
	.emptyEast(emptyProc29East),
	.dataInEast(dataInProc29East),
	.wrEast(wrProc29East),
	.fullEast(fullProc29East),
	.dataOutEast(dataOutProc29East),
	.rdWest(rdProc29West),
	.emptyWest(emptyProc29West),
	.dataInWest(dataInProc29West),
	.wrWest(wrProc29West),
	.fullWest(fullProc29West),
	.dataOutWest(dataOutProc29West));
 
//PROCESSOR 30
system proc30(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe30),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe30),
	.rdNorth(rdProc30North),
	.emptyNorth(emptyProc30North),
	.dataInNorth(dataInProc30North),
	.wrNorth(wrProc30North),
	.fullNorth(fullProc30North),
	.dataOutNorth(dataOutProc30North),
	.rdSouth(rdProc30South),
	.emptySouth(emptyProc30South),
	.dataInSouth(dataInProc30South),
	.wrSouth(wrProc30South),
	.fullSouth(fullProc30South),
	.dataOutSouth(dataOutProc30South),
	.rdEast(rdProc30East),
	.emptyEast(emptyProc30East),
	.dataInEast(dataInProc30East),
	.wrEast(wrProc30East),
	.fullEast(fullProc30East),
	.dataOutEast(dataOutProc30East),
	.rdWest(rdProc30West),
	.emptyWest(emptyProc30West),
	.dataInWest(dataInProc30West),
	.wrWest(wrProc30West),
	.fullWest(fullProc30West),
	.dataOutWest(dataOutProc30West));
 
//PROCESSOR 31
system proc31(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe31),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe31),
	.rdNorth(rdProc31North),
	.emptyNorth(emptyProc31North),
	.dataInNorth(dataInProc31North),
	.wrNorth(wrProc31North),
	.fullNorth(fullProc31North),
	.dataOutNorth(dataOutProc31North),
	.rdSouth(rdProc31South),
	.emptySouth(emptyProc31South),
	.dataInSouth(dataInProc31South),
	.wrSouth(wrProc31South),
	.fullSouth(fullProc31South),
	.dataOutSouth(dataOutProc31South),
	.rdEast(rdProc31East),
	.emptyEast(emptyProc31East),
	.dataInEast(dataInProc31East),
	.wrEast(wrProc31East),
	.fullEast(fullProc31East),
	.dataOutEast(dataOutProc31East),
	.rdWest(rdProc31West),
	.emptyWest(emptyProc31West),
	.dataInWest(dataInProc31West),
	.wrWest(wrProc31West),
	.fullWest(fullProc31West),
	.dataOutWest(dataOutProc31West));
 
//PROCESSOR 32
system proc32(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe32),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe32),
	.rdNorth(rdProc32North),
	.emptyNorth(emptyProc32North),
	.dataInNorth(dataInProc32North),
	.wrNorth(wrProc32North),
	.fullNorth(fullProc32North),
	.dataOutNorth(dataOutProc32North),
	.rdSouth(rdProc32South),
	.emptySouth(emptyProc32South),
	.dataInSouth(dataInProc32South),
	.wrSouth(wrProc32South),
	.fullSouth(fullProc32South),
	.dataOutSouth(dataOutProc32South),
	.rdEast(rdProc32East),
	.emptyEast(emptyProc32East),
	.dataInEast(dataInProc32East),
	.wrEast(wrProc32East),
	.fullEast(fullProc32East),
	.dataOutEast(dataOutProc32East),
	.rdWest(rdProc32West),
	.emptyWest(emptyProc32West),
	.dataInWest(dataInProc32West),
	.wrWest(wrProc32West),
	.fullWest(fullProc32West),
	.dataOutWest(dataOutProc32West));
 
//PROCESSOR 33
system proc33(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe33),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe33),
	.rdNorth(rdProc33North),
	.emptyNorth(emptyProc33North),
	.dataInNorth(dataInProc33North),
	.wrNorth(wrProc33North),
	.fullNorth(fullProc33North),
	.dataOutNorth(dataOutProc33North),
	.rdSouth(rdProc33South),
	.emptySouth(emptyProc33South),
	.dataInSouth(dataInProc33South),
	.wrSouth(wrProc33South),
	.fullSouth(fullProc33South),
	.dataOutSouth(dataOutProc33South),
	.rdEast(rdProc33East),
	.emptyEast(emptyProc33East),
	.dataInEast(dataInProc33East),
	.wrEast(wrProc33East),
	.fullEast(fullProc33East),
	.dataOutEast(dataOutProc33East),
	.rdWest(rdProc33West),
	.emptyWest(emptyProc33West),
	.dataInWest(dataInProc33West),
	.wrWest(wrProc33West),
	.fullWest(fullProc33West),
	.dataOutWest(dataOutProc33West));
 
//PROCESSOR 34
system proc34(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe34),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe34),
	.rdNorth(rdProc34North),
	.emptyNorth(emptyProc34North),
	.dataInNorth(dataInProc34North),
	.wrNorth(wrProc34North),
	.fullNorth(fullProc34North),
	.dataOutNorth(dataOutProc34North),
	.rdSouth(rdProc34South),
	.emptySouth(emptyProc34South),
	.dataInSouth(dataInProc34South),
	.wrSouth(wrProc34South),
	.fullSouth(fullProc34South),
	.dataOutSouth(dataOutProc34South),
	.rdEast(rdProc34East),
	.emptyEast(emptyProc34East),
	.dataInEast(dataInProc34East),
	.wrEast(wrProc34East),
	.fullEast(fullProc34East),
	.dataOutEast(dataOutProc34East),
	.rdWest(rdProc34West),
	.emptyWest(emptyProc34West),
	.dataInWest(dataInProc34West),
	.wrWest(wrProc34West),
	.fullWest(fullProc34West),
	.dataOutWest(dataOutProc34West));
 
//PROCESSOR 35
system proc35(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe35),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe35),
	.rdNorth(rdProc35North),
	.emptyNorth(emptyProc35North),
	.dataInNorth(dataInProc35North),
	.wrNorth(wrProc35North),
	.fullNorth(fullProc35North),
	.dataOutNorth(dataOutProc35North),
	.rdSouth(rdProc35South),
	.emptySouth(emptyProc35South),
	.dataInSouth(dataInProc35South),
	.wrSouth(wrProc35South),
	.fullSouth(fullProc35South),
	.dataOutSouth(dataOutProc35South),
	.rdEast(rdProc35East),
	.emptyEast(emptyProc35East),
	.dataInEast(dataInProc35East),
	.wrEast(wrProc35East),
	.fullEast(fullProc35East),
	.dataOutEast(dataOutProc35East),
	.rdWest(rdProc35West),
	.emptyWest(emptyProc35West),
	.dataInWest(dataInProc35West),
	.wrWest(wrProc35West),
	.fullWest(fullProc35West),
	.dataOutWest(dataOutProc35West));
 
//PROCESSOR 36
system proc36(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe36),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe36),
	.rdNorth(rdProc36North),
	.emptyNorth(emptyProc36North),
	.dataInNorth(dataInProc36North),
	.wrNorth(wrProc36North),
	.fullNorth(fullProc36North),
	.dataOutNorth(dataOutProc36North),
	.rdSouth(rdProc36South),
	.emptySouth(emptyProc36South),
	.dataInSouth(dataInProc36South),
	.wrSouth(wrProc36South),
	.fullSouth(fullProc36South),
	.dataOutSouth(dataOutProc36South),
	.rdEast(rdProc36East),
	.emptyEast(emptyProc36East),
	.dataInEast(dataInProc36East),
	.wrEast(wrProc36East),
	.fullEast(fullProc36East),
	.dataOutEast(dataOutProc36East),
	.rdWest(rdProc36West),
	.emptyWest(emptyProc36West),
	.dataInWest(dataInProc36West),
	.wrWest(wrProc36West),
	.fullWest(fullProc36West),
	.dataOutWest(dataOutProc36West));
 
//PROCESSOR 37
system proc37(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe37),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe37),
	.rdNorth(rdProc37North),
	.emptyNorth(emptyProc37North),
	.dataInNorth(dataInProc37North),
	.wrNorth(wrProc37North),
	.fullNorth(fullProc37North),
	.dataOutNorth(dataOutProc37North),
	.rdSouth(rdProc37South),
	.emptySouth(emptyProc37South),
	.dataInSouth(dataInProc37South),
	.wrSouth(wrProc37South),
	.fullSouth(fullProc37South),
	.dataOutSouth(dataOutProc37South),
	.rdEast(rdProc37East),
	.emptyEast(emptyProc37East),
	.dataInEast(dataInProc37East),
	.wrEast(wrProc37East),
	.fullEast(fullProc37East),
	.dataOutEast(dataOutProc37East),
	.rdWest(rdProc37West),
	.emptyWest(emptyProc37West),
	.dataInWest(dataInProc37West),
	.wrWest(wrProc37West),
	.fullWest(fullProc37West),
	.dataOutWest(dataOutProc37West));
 
//PROCESSOR 38
system proc38(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe38),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe38),
	.rdNorth(rdProc38North),
	.emptyNorth(emptyProc38North),
	.dataInNorth(dataInProc38North),
	.wrNorth(wrProc38North),
	.fullNorth(fullProc38North),
	.dataOutNorth(dataOutProc38North),
	.rdSouth(rdProc38South),
	.emptySouth(emptyProc38South),
	.dataInSouth(dataInProc38South),
	.wrSouth(wrProc38South),
	.fullSouth(fullProc38South),
	.dataOutSouth(dataOutProc38South),
	.rdWest(rdProc38West),
	.emptyWest(emptyProc38West),
	.dataInWest(dataInProc38West),
	.wrWest(wrProc38West),
	.fullWest(fullProc38West),
	.dataOutWest(dataOutProc38West));
 
//PROCESSOR 39
system proc39(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe39),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe39),
	.wrNorth(wrProc39North),
	.fullNorth(fullProc39North),
	.dataOutNorth(dataOutProc39North),
	.rdNorth(rdProc39North),
	.emptyNorth(emptyProc39North),
	.dataInNorth(dataInProc39North),
	.rdSouth(rdProc39South),
	.emptySouth(emptyProc39South),
	.dataInSouth(dataInProc39South),
	.wrSouth(wrProc39South),
	.fullSouth(fullProc39South),
	.dataOutSouth(dataOutProc39South),
	.rdEast(rdProc39East),
	.emptyEast(emptyProc39East),
	.dataInEast(dataInProc39East),
	.wrEast(wrProc39East),
	.fullEast(fullProc39East),
	.dataOutEast(dataOutProc39East));
 
//PROCESSOR 40
system proc40(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe40),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe40),
	.rdNorth(rdProc40North),
	.emptyNorth(emptyProc40North),
	.dataInNorth(dataInProc40North),
	.wrNorth(wrProc40North),
	.fullNorth(fullProc40North),
	.dataOutNorth(dataOutProc40North),
	.rdSouth(rdProc40South),
	.emptySouth(emptyProc40South),
	.dataInSouth(dataInProc40South),
	.wrSouth(wrProc40South),
	.fullSouth(fullProc40South),
	.dataOutSouth(dataOutProc40South),
	.rdEast(rdProc40East),
	.emptyEast(emptyProc40East),
	.dataInEast(dataInProc40East),
	.wrEast(wrProc40East),
	.fullEast(fullProc40East),
	.dataOutEast(dataOutProc40East),
	.rdWest(rdProc40West),
	.emptyWest(emptyProc40West),
	.dataInWest(dataInProc40West),
	.wrWest(wrProc40West),
	.fullWest(fullProc40West),
	.dataOutWest(dataOutProc40West));
 
//PROCESSOR 41
system proc41(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe41),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe41),
	.rdNorth(rdProc41North),
	.emptyNorth(emptyProc41North),
	.dataInNorth(dataInProc41North),
	.wrNorth(wrProc41North),
	.fullNorth(fullProc41North),
	.dataOutNorth(dataOutProc41North),
	.rdSouth(rdProc41South),
	.emptySouth(emptyProc41South),
	.dataInSouth(dataInProc41South),
	.wrSouth(wrProc41South),
	.fullSouth(fullProc41South),
	.dataOutSouth(dataOutProc41South),
	.rdEast(rdProc41East),
	.emptyEast(emptyProc41East),
	.dataInEast(dataInProc41East),
	.wrEast(wrProc41East),
	.fullEast(fullProc41East),
	.dataOutEast(dataOutProc41East),
	.rdWest(rdProc41West),
	.emptyWest(emptyProc41West),
	.dataInWest(dataInProc41West),
	.wrWest(wrProc41West),
	.fullWest(fullProc41West),
	.dataOutWest(dataOutProc41West));
 
//PROCESSOR 42
system proc42(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe42),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe42),
	.rdNorth(rdProc42North),
	.emptyNorth(emptyProc42North),
	.dataInNorth(dataInProc42North),
	.wrNorth(wrProc42North),
	.fullNorth(fullProc42North),
	.dataOutNorth(dataOutProc42North),
	.rdSouth(rdProc42South),
	.emptySouth(emptyProc42South),
	.dataInSouth(dataInProc42South),
	.wrSouth(wrProc42South),
	.fullSouth(fullProc42South),
	.dataOutSouth(dataOutProc42South),
	.rdEast(rdProc42East),
	.emptyEast(emptyProc42East),
	.dataInEast(dataInProc42East),
	.wrEast(wrProc42East),
	.fullEast(fullProc42East),
	.dataOutEast(dataOutProc42East),
	.rdWest(rdProc42West),
	.emptyWest(emptyProc42West),
	.dataInWest(dataInProc42West),
	.wrWest(wrProc42West),
	.fullWest(fullProc42West),
	.dataOutWest(dataOutProc42West));
 
//PROCESSOR 43
system proc43(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe43),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe43),
	.rdNorth(rdProc43North),
	.emptyNorth(emptyProc43North),
	.dataInNorth(dataInProc43North),
	.wrNorth(wrProc43North),
	.fullNorth(fullProc43North),
	.dataOutNorth(dataOutProc43North),
	.rdSouth(rdProc43South),
	.emptySouth(emptyProc43South),
	.dataInSouth(dataInProc43South),
	.wrSouth(wrProc43South),
	.fullSouth(fullProc43South),
	.dataOutSouth(dataOutProc43South),
	.rdEast(rdProc43East),
	.emptyEast(emptyProc43East),
	.dataInEast(dataInProc43East),
	.wrEast(wrProc43East),
	.fullEast(fullProc43East),
	.dataOutEast(dataOutProc43East),
	.rdWest(rdProc43West),
	.emptyWest(emptyProc43West),
	.dataInWest(dataInProc43West),
	.wrWest(wrProc43West),
	.fullWest(fullProc43West),
	.dataOutWest(dataOutProc43West));
 
//PROCESSOR 44
system proc44(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe44),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe44),
	.rdNorth(rdProc44North),
	.emptyNorth(emptyProc44North),
	.dataInNorth(dataInProc44North),
	.wrNorth(wrProc44North),
	.fullNorth(fullProc44North),
	.dataOutNorth(dataOutProc44North),
	.rdSouth(rdProc44South),
	.emptySouth(emptyProc44South),
	.dataInSouth(dataInProc44South),
	.wrSouth(wrProc44South),
	.fullSouth(fullProc44South),
	.dataOutSouth(dataOutProc44South),
	.rdEast(rdProc44East),
	.emptyEast(emptyProc44East),
	.dataInEast(dataInProc44East),
	.wrEast(wrProc44East),
	.fullEast(fullProc44East),
	.dataOutEast(dataOutProc44East),
	.rdWest(rdProc44West),
	.emptyWest(emptyProc44West),
	.dataInWest(dataInProc44West),
	.wrWest(wrProc44West),
	.fullWest(fullProc44West),
	.dataOutWest(dataOutProc44West));
 
//PROCESSOR 45
system proc45(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe45),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe45),
	.rdNorth(rdProc45North),
	.emptyNorth(emptyProc45North),
	.dataInNorth(dataInProc45North),
	.wrNorth(wrProc45North),
	.fullNorth(fullProc45North),
	.dataOutNorth(dataOutProc45North),
	.rdSouth(rdProc45South),
	.emptySouth(emptyProc45South),
	.dataInSouth(dataInProc45South),
	.wrSouth(wrProc45South),
	.fullSouth(fullProc45South),
	.dataOutSouth(dataOutProc45South),
	.rdEast(rdProc45East),
	.emptyEast(emptyProc45East),
	.dataInEast(dataInProc45East),
	.wrEast(wrProc45East),
	.fullEast(fullProc45East),
	.dataOutEast(dataOutProc45East),
	.rdWest(rdProc45West),
	.emptyWest(emptyProc45West),
	.dataInWest(dataInProc45West),
	.wrWest(wrProc45West),
	.fullWest(fullProc45West),
	.dataOutWest(dataOutProc45West));
 
//PROCESSOR 46
system proc46(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe46),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe46),
	.rdNorth(rdProc46North),
	.emptyNorth(emptyProc46North),
	.dataInNorth(dataInProc46North),
	.wrNorth(wrProc46North),
	.fullNorth(fullProc46North),
	.dataOutNorth(dataOutProc46North),
	.rdSouth(rdProc46South),
	.emptySouth(emptyProc46South),
	.dataInSouth(dataInProc46South),
	.wrSouth(wrProc46South),
	.fullSouth(fullProc46South),
	.dataOutSouth(dataOutProc46South),
	.rdEast(rdProc46East),
	.emptyEast(emptyProc46East),
	.dataInEast(dataInProc46East),
	.wrEast(wrProc46East),
	.fullEast(fullProc46East),
	.dataOutEast(dataOutProc46East),
	.rdWest(rdProc46West),
	.emptyWest(emptyProc46West),
	.dataInWest(dataInProc46West),
	.wrWest(wrProc46West),
	.fullWest(fullProc46West),
	.dataOutWest(dataOutProc46West));
 
//PROCESSOR 47
system proc47(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe47),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe47),
	.rdNorth(rdProc47North),
	.emptyNorth(emptyProc47North),
	.dataInNorth(dataInProc47North),
	.wrNorth(wrProc47North),
	.fullNorth(fullProc47North),
	.dataOutNorth(dataOutProc47North),
	.rdSouth(rdProc47South),
	.emptySouth(emptyProc47South),
	.dataInSouth(dataInProc47South),
	.wrSouth(wrProc47South),
	.fullSouth(fullProc47South),
	.dataOutSouth(dataOutProc47South),
	.rdEast(rdProc47East),
	.emptyEast(emptyProc47East),
	.dataInEast(dataInProc47East),
	.wrEast(wrProc47East),
	.fullEast(fullProc47East),
	.dataOutEast(dataOutProc47East),
	.rdWest(rdProc47West),
	.emptyWest(emptyProc47West),
	.dataInWest(dataInProc47West),
	.wrWest(wrProc47West),
	.fullWest(fullProc47West),
	.dataOutWest(dataOutProc47West));
 
//PROCESSOR 48
system proc48(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe48),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe48),
	.rdNorth(rdProc48North),
	.emptyNorth(emptyProc48North),
	.dataInNorth(dataInProc48North),
	.wrNorth(wrProc48North),
	.fullNorth(fullProc48North),
	.dataOutNorth(dataOutProc48North),
	.rdSouth(rdProc48South),
	.emptySouth(emptyProc48South),
	.dataInSouth(dataInProc48South),
	.wrSouth(wrProc48South),
	.fullSouth(fullProc48South),
	.dataOutSouth(dataOutProc48South),
	.rdEast(rdProc48East),
	.emptyEast(emptyProc48East),
	.dataInEast(dataInProc48East),
	.wrEast(wrProc48East),
	.fullEast(fullProc48East),
	.dataOutEast(dataOutProc48East),
	.rdWest(rdProc48West),
	.emptyWest(emptyProc48West),
	.dataInWest(dataInProc48West),
	.wrWest(wrProc48West),
	.fullWest(fullProc48West),
	.dataOutWest(dataOutProc48West));
 
//PROCESSOR 49
system proc49(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe49),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe49),
	.rdNorth(rdProc49North),
	.emptyNorth(emptyProc49North),
	.dataInNorth(dataInProc49North),
	.wrNorth(wrProc49North),
	.fullNorth(fullProc49North),
	.dataOutNorth(dataOutProc49North),
	.rdSouth(rdProc49South),
	.emptySouth(emptyProc49South),
	.dataInSouth(dataInProc49South),
	.wrSouth(wrProc49South),
	.fullSouth(fullProc49South),
	.dataOutSouth(dataOutProc49South),
	.rdEast(rdProc49East),
	.emptyEast(emptyProc49East),
	.dataInEast(dataInProc49East),
	.wrEast(wrProc49East),
	.fullEast(fullProc49East),
	.dataOutEast(dataOutProc49East),
	.rdWest(rdProc49West),
	.emptyWest(emptyProc49West),
	.dataInWest(dataInProc49West),
	.wrWest(wrProc49West),
	.fullWest(fullProc49West),
	.dataOutWest(dataOutProc49West));
 
//PROCESSOR 50
system proc50(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe50),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe50),
	.rdNorth(rdProc50North),
	.emptyNorth(emptyProc50North),
	.dataInNorth(dataInProc50North),
	.wrNorth(wrProc50North),
	.fullNorth(fullProc50North),
	.dataOutNorth(dataOutProc50North),
	.rdSouth(rdProc50South),
	.emptySouth(emptyProc50South),
	.dataInSouth(dataInProc50South),
	.wrSouth(wrProc50South),
	.fullSouth(fullProc50South),
	.dataOutSouth(dataOutProc50South),
	.rdEast(rdProc50East),
	.emptyEast(emptyProc50East),
	.dataInEast(dataInProc50East),
	.wrEast(wrProc50East),
	.fullEast(fullProc50East),
	.dataOutEast(dataOutProc50East),
	.rdWest(rdProc50West),
	.emptyWest(emptyProc50West),
	.dataInWest(dataInProc50West),
	.wrWest(wrProc50West),
	.fullWest(fullProc50West),
	.dataOutWest(dataOutProc50West));
 
//PROCESSOR 51
system proc51(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe51),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe51),
	.rdNorth(rdProc51North),
	.emptyNorth(emptyProc51North),
	.dataInNorth(dataInProc51North),
	.wrNorth(wrProc51North),
	.fullNorth(fullProc51North),
	.dataOutNorth(dataOutProc51North),
	.rdSouth(rdProc51South),
	.emptySouth(emptyProc51South),
	.dataInSouth(dataInProc51South),
	.wrSouth(wrProc51South),
	.fullSouth(fullProc51South),
	.dataOutSouth(dataOutProc51South),
	.rdWest(rdProc51West),
	.emptyWest(emptyProc51West),
	.dataInWest(dataInProc51West),
	.wrWest(wrProc51West),
	.fullWest(fullProc51West),
	.dataOutWest(dataOutProc51West));
 
//PROCESSOR 52
system proc52(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe52),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe52),
	.wrNorth(wrProc52North),
	.fullNorth(fullProc52North),
	.dataOutNorth(dataOutProc52North),
	.rdNorth(rdProc52North),
	.emptyNorth(emptyProc52North),
	.dataInNorth(dataInProc52North),
	.rdSouth(rdProc52South),
	.emptySouth(emptyProc52South),
	.dataInSouth(dataInProc52South),
	.wrSouth(wrProc52South),
	.fullSouth(fullProc52South),
	.dataOutSouth(dataOutProc52South),
	.rdEast(rdProc52East),
	.emptyEast(emptyProc52East),
	.dataInEast(dataInProc52East),
	.wrEast(wrProc52East),
	.fullEast(fullProc52East),
	.dataOutEast(dataOutProc52East));
 
//PROCESSOR 53
system proc53(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe53),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe53),
	.rdNorth(rdProc53North),
	.emptyNorth(emptyProc53North),
	.dataInNorth(dataInProc53North),
	.wrNorth(wrProc53North),
	.fullNorth(fullProc53North),
	.dataOutNorth(dataOutProc53North),
	.rdSouth(rdProc53South),
	.emptySouth(emptyProc53South),
	.dataInSouth(dataInProc53South),
	.wrSouth(wrProc53South),
	.fullSouth(fullProc53South),
	.dataOutSouth(dataOutProc53South),
	.rdEast(rdProc53East),
	.emptyEast(emptyProc53East),
	.dataInEast(dataInProc53East),
	.wrEast(wrProc53East),
	.fullEast(fullProc53East),
	.dataOutEast(dataOutProc53East),
	.rdWest(rdProc53West),
	.emptyWest(emptyProc53West),
	.dataInWest(dataInProc53West),
	.wrWest(wrProc53West),
	.fullWest(fullProc53West),
	.dataOutWest(dataOutProc53West));
 
//PROCESSOR 54
system proc54(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe54),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe54),
	.rdNorth(rdProc54North),
	.emptyNorth(emptyProc54North),
	.dataInNorth(dataInProc54North),
	.wrNorth(wrProc54North),
	.fullNorth(fullProc54North),
	.dataOutNorth(dataOutProc54North),
	.rdSouth(rdProc54South),
	.emptySouth(emptyProc54South),
	.dataInSouth(dataInProc54South),
	.wrSouth(wrProc54South),
	.fullSouth(fullProc54South),
	.dataOutSouth(dataOutProc54South),
	.rdEast(rdProc54East),
	.emptyEast(emptyProc54East),
	.dataInEast(dataInProc54East),
	.wrEast(wrProc54East),
	.fullEast(fullProc54East),
	.dataOutEast(dataOutProc54East),
	.rdWest(rdProc54West),
	.emptyWest(emptyProc54West),
	.dataInWest(dataInProc54West),
	.wrWest(wrProc54West),
	.fullWest(fullProc54West),
	.dataOutWest(dataOutProc54West));
 
//PROCESSOR 55
system proc55(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe55),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe55),
	.rdNorth(rdProc55North),
	.emptyNorth(emptyProc55North),
	.dataInNorth(dataInProc55North),
	.wrNorth(wrProc55North),
	.fullNorth(fullProc55North),
	.dataOutNorth(dataOutProc55North),
	.rdSouth(rdProc55South),
	.emptySouth(emptyProc55South),
	.dataInSouth(dataInProc55South),
	.wrSouth(wrProc55South),
	.fullSouth(fullProc55South),
	.dataOutSouth(dataOutProc55South),
	.rdEast(rdProc55East),
	.emptyEast(emptyProc55East),
	.dataInEast(dataInProc55East),
	.wrEast(wrProc55East),
	.fullEast(fullProc55East),
	.dataOutEast(dataOutProc55East),
	.rdWest(rdProc55West),
	.emptyWest(emptyProc55West),
	.dataInWest(dataInProc55West),
	.wrWest(wrProc55West),
	.fullWest(fullProc55West),
	.dataOutWest(dataOutProc55West));
 
//PROCESSOR 56
system proc56(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe56),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe56),
	.rdNorth(rdProc56North),
	.emptyNorth(emptyProc56North),
	.dataInNorth(dataInProc56North),
	.wrNorth(wrProc56North),
	.fullNorth(fullProc56North),
	.dataOutNorth(dataOutProc56North),
	.rdSouth(rdProc56South),
	.emptySouth(emptyProc56South),
	.dataInSouth(dataInProc56South),
	.wrSouth(wrProc56South),
	.fullSouth(fullProc56South),
	.dataOutSouth(dataOutProc56South),
	.rdEast(rdProc56East),
	.emptyEast(emptyProc56East),
	.dataInEast(dataInProc56East),
	.wrEast(wrProc56East),
	.fullEast(fullProc56East),
	.dataOutEast(dataOutProc56East),
	.rdWest(rdProc56West),
	.emptyWest(emptyProc56West),
	.dataInWest(dataInProc56West),
	.wrWest(wrProc56West),
	.fullWest(fullProc56West),
	.dataOutWest(dataOutProc56West));
 
//PROCESSOR 57
system proc57(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe57),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe57),
	.rdNorth(rdProc57North),
	.emptyNorth(emptyProc57North),
	.dataInNorth(dataInProc57North),
	.wrNorth(wrProc57North),
	.fullNorth(fullProc57North),
	.dataOutNorth(dataOutProc57North),
	.rdSouth(rdProc57South),
	.emptySouth(emptyProc57South),
	.dataInSouth(dataInProc57South),
	.wrSouth(wrProc57South),
	.fullSouth(fullProc57South),
	.dataOutSouth(dataOutProc57South),
	.rdEast(rdProc57East),
	.emptyEast(emptyProc57East),
	.dataInEast(dataInProc57East),
	.wrEast(wrProc57East),
	.fullEast(fullProc57East),
	.dataOutEast(dataOutProc57East),
	.rdWest(rdProc57West),
	.emptyWest(emptyProc57West),
	.dataInWest(dataInProc57West),
	.wrWest(wrProc57West),
	.fullWest(fullProc57West),
	.dataOutWest(dataOutProc57West));
 
//PROCESSOR 58
system proc58(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe58),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe58),
	.rdNorth(rdProc58North),
	.emptyNorth(emptyProc58North),
	.dataInNorth(dataInProc58North),
	.wrNorth(wrProc58North),
	.fullNorth(fullProc58North),
	.dataOutNorth(dataOutProc58North),
	.rdSouth(rdProc58South),
	.emptySouth(emptyProc58South),
	.dataInSouth(dataInProc58South),
	.wrSouth(wrProc58South),
	.fullSouth(fullProc58South),
	.dataOutSouth(dataOutProc58South),
	.rdEast(rdProc58East),
	.emptyEast(emptyProc58East),
	.dataInEast(dataInProc58East),
	.wrEast(wrProc58East),
	.fullEast(fullProc58East),
	.dataOutEast(dataOutProc58East),
	.rdWest(rdProc58West),
	.emptyWest(emptyProc58West),
	.dataInWest(dataInProc58West),
	.wrWest(wrProc58West),
	.fullWest(fullProc58West),
	.dataOutWest(dataOutProc58West));
 
//PROCESSOR 59
system proc59(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe59),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe59),
	.rdNorth(rdProc59North),
	.emptyNorth(emptyProc59North),
	.dataInNorth(dataInProc59North),
	.wrNorth(wrProc59North),
	.fullNorth(fullProc59North),
	.dataOutNorth(dataOutProc59North),
	.rdSouth(rdProc59South),
	.emptySouth(emptyProc59South),
	.dataInSouth(dataInProc59South),
	.wrSouth(wrProc59South),
	.fullSouth(fullProc59South),
	.dataOutSouth(dataOutProc59South),
	.rdEast(rdProc59East),
	.emptyEast(emptyProc59East),
	.dataInEast(dataInProc59East),
	.wrEast(wrProc59East),
	.fullEast(fullProc59East),
	.dataOutEast(dataOutProc59East),
	.rdWest(rdProc59West),
	.emptyWest(emptyProc59West),
	.dataInWest(dataInProc59West),
	.wrWest(wrProc59West),
	.fullWest(fullProc59West),
	.dataOutWest(dataOutProc59West));
 
//PROCESSOR 60
system proc60(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe60),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe60),
	.rdNorth(rdProc60North),
	.emptyNorth(emptyProc60North),
	.dataInNorth(dataInProc60North),
	.wrNorth(wrProc60North),
	.fullNorth(fullProc60North),
	.dataOutNorth(dataOutProc60North),
	.rdSouth(rdProc60South),
	.emptySouth(emptyProc60South),
	.dataInSouth(dataInProc60South),
	.wrSouth(wrProc60South),
	.fullSouth(fullProc60South),
	.dataOutSouth(dataOutProc60South),
	.rdEast(rdProc60East),
	.emptyEast(emptyProc60East),
	.dataInEast(dataInProc60East),
	.wrEast(wrProc60East),
	.fullEast(fullProc60East),
	.dataOutEast(dataOutProc60East),
	.rdWest(rdProc60West),
	.emptyWest(emptyProc60West),
	.dataInWest(dataInProc60West),
	.wrWest(wrProc60West),
	.fullWest(fullProc60West),
	.dataOutWest(dataOutProc60West));
 
//PROCESSOR 61
system proc61(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe61),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe61),
	.rdNorth(rdProc61North),
	.emptyNorth(emptyProc61North),
	.dataInNorth(dataInProc61North),
	.wrNorth(wrProc61North),
	.fullNorth(fullProc61North),
	.dataOutNorth(dataOutProc61North),
	.rdSouth(rdProc61South),
	.emptySouth(emptyProc61South),
	.dataInSouth(dataInProc61South),
	.wrSouth(wrProc61South),
	.fullSouth(fullProc61South),
	.dataOutSouth(dataOutProc61South),
	.rdEast(rdProc61East),
	.emptyEast(emptyProc61East),
	.dataInEast(dataInProc61East),
	.wrEast(wrProc61East),
	.fullEast(fullProc61East),
	.dataOutEast(dataOutProc61East),
	.rdWest(rdProc61West),
	.emptyWest(emptyProc61West),
	.dataInWest(dataInProc61West),
	.wrWest(wrProc61West),
	.fullWest(fullProc61West),
	.dataOutWest(dataOutProc61West));
 
//PROCESSOR 62
system proc62(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe62),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe62),
	.rdNorth(rdProc62North),
	.emptyNorth(emptyProc62North),
	.dataInNorth(dataInProc62North),
	.wrNorth(wrProc62North),
	.fullNorth(fullProc62North),
	.dataOutNorth(dataOutProc62North),
	.rdSouth(rdProc62South),
	.emptySouth(emptyProc62South),
	.dataInSouth(dataInProc62South),
	.wrSouth(wrProc62South),
	.fullSouth(fullProc62South),
	.dataOutSouth(dataOutProc62South),
	.rdEast(rdProc62East),
	.emptyEast(emptyProc62East),
	.dataInEast(dataInProc62East),
	.wrEast(wrProc62East),
	.fullEast(fullProc62East),
	.dataOutEast(dataOutProc62East),
	.rdWest(rdProc62West),
	.emptyWest(emptyProc62West),
	.dataInWest(dataInProc62West),
	.wrWest(wrProc62West),
	.fullWest(fullProc62West),
	.dataOutWest(dataOutProc62West));
 
//PROCESSOR 63
system proc63(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe63),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe63),
	.rdNorth(rdProc63North),
	.emptyNorth(emptyProc63North),
	.dataInNorth(dataInProc63North),
	.wrNorth(wrProc63North),
	.fullNorth(fullProc63North),
	.dataOutNorth(dataOutProc63North),
	.rdSouth(rdProc63South),
	.emptySouth(emptyProc63South),
	.dataInSouth(dataInProc63South),
	.wrSouth(wrProc63South),
	.fullSouth(fullProc63South),
	.dataOutSouth(dataOutProc63South),
	.rdEast(rdProc63East),
	.emptyEast(emptyProc63East),
	.dataInEast(dataInProc63East),
	.wrEast(wrProc63East),
	.fullEast(fullProc63East),
	.dataOutEast(dataOutProc63East),
	.rdWest(rdProc63West),
	.emptyWest(emptyProc63West),
	.dataInWest(dataInProc63West),
	.wrWest(wrProc63West),
	.fullWest(fullProc63West),
	.dataOutWest(dataOutProc63West));
 
//PROCESSOR 64
system proc64(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe64),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe64),
	.rdNorth(rdProc64North),
	.emptyNorth(emptyProc64North),
	.dataInNorth(dataInProc64North),
	.wrNorth(wrProc64North),
	.fullNorth(fullProc64North),
	.dataOutNorth(dataOutProc64North),
	.rdSouth(rdProc64South),
	.emptySouth(emptyProc64South),
	.dataInSouth(dataInProc64South),
	.wrSouth(wrProc64South),
	.fullSouth(fullProc64South),
	.dataOutSouth(dataOutProc64South),
	.rdWest(rdProc64West),
	.emptyWest(emptyProc64West),
	.dataInWest(dataInProc64West),
	.wrWest(wrProc64West),
	.fullWest(fullProc64West),
	.dataOutWest(dataOutProc64West));
 
//PROCESSOR 65
system proc65(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe65),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe65),
	.wrNorth(wrProc65North),
	.fullNorth(fullProc65North),
	.dataOutNorth(dataOutProc65North),
	.rdNorth(rdProc65North),
	.emptyNorth(emptyProc65North),
	.dataInNorth(dataInProc65North),
	.rdSouth(rdProc65South),
	.emptySouth(emptyProc65South),
	.dataInSouth(dataInProc65South),
	.wrSouth(wrProc65South),
	.fullSouth(fullProc65South),
	.dataOutSouth(dataOutProc65South),
	.rdEast(rdProc65East),
	.emptyEast(emptyProc65East),
	.dataInEast(dataInProc65East),
	.wrEast(wrProc65East),
	.fullEast(fullProc65East),
	.dataOutEast(dataOutProc65East));
 
//PROCESSOR 66
system proc66(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe66),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe66),
	.rdNorth(rdProc66North),
	.emptyNorth(emptyProc66North),
	.dataInNorth(dataInProc66North),
	.wrNorth(wrProc66North),
	.fullNorth(fullProc66North),
	.dataOutNorth(dataOutProc66North),
	.rdSouth(rdProc66South),
	.emptySouth(emptyProc66South),
	.dataInSouth(dataInProc66South),
	.wrSouth(wrProc66South),
	.fullSouth(fullProc66South),
	.dataOutSouth(dataOutProc66South),
	.rdEast(rdProc66East),
	.emptyEast(emptyProc66East),
	.dataInEast(dataInProc66East),
	.wrEast(wrProc66East),
	.fullEast(fullProc66East),
	.dataOutEast(dataOutProc66East),
	.rdWest(rdProc66West),
	.emptyWest(emptyProc66West),
	.dataInWest(dataInProc66West),
	.wrWest(wrProc66West),
	.fullWest(fullProc66West),
	.dataOutWest(dataOutProc66West));
 
//PROCESSOR 67
system proc67(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe67),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe67),
	.rdNorth(rdProc67North),
	.emptyNorth(emptyProc67North),
	.dataInNorth(dataInProc67North),
	.wrNorth(wrProc67North),
	.fullNorth(fullProc67North),
	.dataOutNorth(dataOutProc67North),
	.rdSouth(rdProc67South),
	.emptySouth(emptyProc67South),
	.dataInSouth(dataInProc67South),
	.wrSouth(wrProc67South),
	.fullSouth(fullProc67South),
	.dataOutSouth(dataOutProc67South),
	.rdEast(rdProc67East),
	.emptyEast(emptyProc67East),
	.dataInEast(dataInProc67East),
	.wrEast(wrProc67East),
	.fullEast(fullProc67East),
	.dataOutEast(dataOutProc67East),
	.rdWest(rdProc67West),
	.emptyWest(emptyProc67West),
	.dataInWest(dataInProc67West),
	.wrWest(wrProc67West),
	.fullWest(fullProc67West),
	.dataOutWest(dataOutProc67West));
 
//PROCESSOR 68
system proc68(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe68),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe68),
	.rdNorth(rdProc68North),
	.emptyNorth(emptyProc68North),
	.dataInNorth(dataInProc68North),
	.wrNorth(wrProc68North),
	.fullNorth(fullProc68North),
	.dataOutNorth(dataOutProc68North),
	.rdSouth(rdProc68South),
	.emptySouth(emptyProc68South),
	.dataInSouth(dataInProc68South),
	.wrSouth(wrProc68South),
	.fullSouth(fullProc68South),
	.dataOutSouth(dataOutProc68South),
	.rdEast(rdProc68East),
	.emptyEast(emptyProc68East),
	.dataInEast(dataInProc68East),
	.wrEast(wrProc68East),
	.fullEast(fullProc68East),
	.dataOutEast(dataOutProc68East),
	.rdWest(rdProc68West),
	.emptyWest(emptyProc68West),
	.dataInWest(dataInProc68West),
	.wrWest(wrProc68West),
	.fullWest(fullProc68West),
	.dataOutWest(dataOutProc68West));
 
//PROCESSOR 69
system proc69(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe69),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe69),
	.rdNorth(rdProc69North),
	.emptyNorth(emptyProc69North),
	.dataInNorth(dataInProc69North),
	.wrNorth(wrProc69North),
	.fullNorth(fullProc69North),
	.dataOutNorth(dataOutProc69North),
	.rdSouth(rdProc69South),
	.emptySouth(emptyProc69South),
	.dataInSouth(dataInProc69South),
	.wrSouth(wrProc69South),
	.fullSouth(fullProc69South),
	.dataOutSouth(dataOutProc69South),
	.rdEast(rdProc69East),
	.emptyEast(emptyProc69East),
	.dataInEast(dataInProc69East),
	.wrEast(wrProc69East),
	.fullEast(fullProc69East),
	.dataOutEast(dataOutProc69East),
	.rdWest(rdProc69West),
	.emptyWest(emptyProc69West),
	.dataInWest(dataInProc69West),
	.wrWest(wrProc69West),
	.fullWest(fullProc69West),
	.dataOutWest(dataOutProc69West));
 
//PROCESSOR 70
system proc70(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe70),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe70),
	.rdNorth(rdProc70North),
	.emptyNorth(emptyProc70North),
	.dataInNorth(dataInProc70North),
	.wrNorth(wrProc70North),
	.fullNorth(fullProc70North),
	.dataOutNorth(dataOutProc70North),
	.rdSouth(rdProc70South),
	.emptySouth(emptyProc70South),
	.dataInSouth(dataInProc70South),
	.wrSouth(wrProc70South),
	.fullSouth(fullProc70South),
	.dataOutSouth(dataOutProc70South),
	.rdEast(rdProc70East),
	.emptyEast(emptyProc70East),
	.dataInEast(dataInProc70East),
	.wrEast(wrProc70East),
	.fullEast(fullProc70East),
	.dataOutEast(dataOutProc70East),
	.rdWest(rdProc70West),
	.emptyWest(emptyProc70West),
	.dataInWest(dataInProc70West),
	.wrWest(wrProc70West),
	.fullWest(fullProc70West),
	.dataOutWest(dataOutProc70West));
 
//PROCESSOR 71
system proc71(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe71),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe71),
	.rdNorth(rdProc71North),
	.emptyNorth(emptyProc71North),
	.dataInNorth(dataInProc71North),
	.wrNorth(wrProc71North),
	.fullNorth(fullProc71North),
	.dataOutNorth(dataOutProc71North),
	.rdSouth(rdProc71South),
	.emptySouth(emptyProc71South),
	.dataInSouth(dataInProc71South),
	.wrSouth(wrProc71South),
	.fullSouth(fullProc71South),
	.dataOutSouth(dataOutProc71South),
	.rdEast(rdProc71East),
	.emptyEast(emptyProc71East),
	.dataInEast(dataInProc71East),
	.wrEast(wrProc71East),
	.fullEast(fullProc71East),
	.dataOutEast(dataOutProc71East),
	.rdWest(rdProc71West),
	.emptyWest(emptyProc71West),
	.dataInWest(dataInProc71West),
	.wrWest(wrProc71West),
	.fullWest(fullProc71West),
	.dataOutWest(dataOutProc71West));
 
//PROCESSOR 72
system proc72(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe72),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe72),
	.rdNorth(rdProc72North),
	.emptyNorth(emptyProc72North),
	.dataInNorth(dataInProc72North),
	.wrNorth(wrProc72North),
	.fullNorth(fullProc72North),
	.dataOutNorth(dataOutProc72North),
	.rdSouth(rdProc72South),
	.emptySouth(emptyProc72South),
	.dataInSouth(dataInProc72South),
	.wrSouth(wrProc72South),
	.fullSouth(fullProc72South),
	.dataOutSouth(dataOutProc72South),
	.rdEast(rdProc72East),
	.emptyEast(emptyProc72East),
	.dataInEast(dataInProc72East),
	.wrEast(wrProc72East),
	.fullEast(fullProc72East),
	.dataOutEast(dataOutProc72East),
	.rdWest(rdProc72West),
	.emptyWest(emptyProc72West),
	.dataInWest(dataInProc72West),
	.wrWest(wrProc72West),
	.fullWest(fullProc72West),
	.dataOutWest(dataOutProc72West));
 
//PROCESSOR 73
system proc73(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe73),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe73),
	.rdNorth(rdProc73North),
	.emptyNorth(emptyProc73North),
	.dataInNorth(dataInProc73North),
	.wrNorth(wrProc73North),
	.fullNorth(fullProc73North),
	.dataOutNorth(dataOutProc73North),
	.rdSouth(rdProc73South),
	.emptySouth(emptyProc73South),
	.dataInSouth(dataInProc73South),
	.wrSouth(wrProc73South),
	.fullSouth(fullProc73South),
	.dataOutSouth(dataOutProc73South),
	.rdEast(rdProc73East),
	.emptyEast(emptyProc73East),
	.dataInEast(dataInProc73East),
	.wrEast(wrProc73East),
	.fullEast(fullProc73East),
	.dataOutEast(dataOutProc73East),
	.rdWest(rdProc73West),
	.emptyWest(emptyProc73West),
	.dataInWest(dataInProc73West),
	.wrWest(wrProc73West),
	.fullWest(fullProc73West),
	.dataOutWest(dataOutProc73West));
 
//PROCESSOR 74
system proc74(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe74),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe74),
	.rdNorth(rdProc74North),
	.emptyNorth(emptyProc74North),
	.dataInNorth(dataInProc74North),
	.wrNorth(wrProc74North),
	.fullNorth(fullProc74North),
	.dataOutNorth(dataOutProc74North),
	.rdSouth(rdProc74South),
	.emptySouth(emptyProc74South),
	.dataInSouth(dataInProc74South),
	.wrSouth(wrProc74South),
	.fullSouth(fullProc74South),
	.dataOutSouth(dataOutProc74South),
	.rdEast(rdProc74East),
	.emptyEast(emptyProc74East),
	.dataInEast(dataInProc74East),
	.wrEast(wrProc74East),
	.fullEast(fullProc74East),
	.dataOutEast(dataOutProc74East),
	.rdWest(rdProc74West),
	.emptyWest(emptyProc74West),
	.dataInWest(dataInProc74West),
	.wrWest(wrProc74West),
	.fullWest(fullProc74West),
	.dataOutWest(dataOutProc74West));
 
//PROCESSOR 75
system proc75(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe75),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe75),
	.rdNorth(rdProc75North),
	.emptyNorth(emptyProc75North),
	.dataInNorth(dataInProc75North),
	.wrNorth(wrProc75North),
	.fullNorth(fullProc75North),
	.dataOutNorth(dataOutProc75North),
	.rdSouth(rdProc75South),
	.emptySouth(emptyProc75South),
	.dataInSouth(dataInProc75South),
	.wrSouth(wrProc75South),
	.fullSouth(fullProc75South),
	.dataOutSouth(dataOutProc75South),
	.rdEast(rdProc75East),
	.emptyEast(emptyProc75East),
	.dataInEast(dataInProc75East),
	.wrEast(wrProc75East),
	.fullEast(fullProc75East),
	.dataOutEast(dataOutProc75East),
	.rdWest(rdProc75West),
	.emptyWest(emptyProc75West),
	.dataInWest(dataInProc75West),
	.wrWest(wrProc75West),
	.fullWest(fullProc75West),
	.dataOutWest(dataOutProc75West));
 
//PROCESSOR 76
system proc76(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe76),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe76),
	.rdNorth(rdProc76North),
	.emptyNorth(emptyProc76North),
	.dataInNorth(dataInProc76North),
	.wrNorth(wrProc76North),
	.fullNorth(fullProc76North),
	.dataOutNorth(dataOutProc76North),
	.rdSouth(rdProc76South),
	.emptySouth(emptyProc76South),
	.dataInSouth(dataInProc76South),
	.wrSouth(wrProc76South),
	.fullSouth(fullProc76South),
	.dataOutSouth(dataOutProc76South),
	.rdEast(rdProc76East),
	.emptyEast(emptyProc76East),
	.dataInEast(dataInProc76East),
	.wrEast(wrProc76East),
	.fullEast(fullProc76East),
	.dataOutEast(dataOutProc76East),
	.rdWest(rdProc76West),
	.emptyWest(emptyProc76West),
	.dataInWest(dataInProc76West),
	.wrWest(wrProc76West),
	.fullWest(fullProc76West),
	.dataOutWest(dataOutProc76West));
 
//PROCESSOR 77
system proc77(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe77),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe77),
	.rdNorth(rdProc77North),
	.emptyNorth(emptyProc77North),
	.dataInNorth(dataInProc77North),
	.wrNorth(wrProc77North),
	.fullNorth(fullProc77North),
	.dataOutNorth(dataOutProc77North),
	.rdSouth(rdProc77South),
	.emptySouth(emptyProc77South),
	.dataInSouth(dataInProc77South),
	.wrSouth(wrProc77South),
	.fullSouth(fullProc77South),
	.dataOutSouth(dataOutProc77South),
	.rdWest(rdProc77West),
	.emptyWest(emptyProc77West),
	.dataInWest(dataInProc77West),
	.wrWest(wrProc77West),
	.fullWest(fullProc77West),
	.dataOutWest(dataOutProc77West));
 
//PROCESSOR 78
system proc78(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe78),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe78),
	.wrNorth(wrProc78North),
	.fullNorth(fullProc78North),
	.dataOutNorth(dataOutProc78North),
	.rdNorth(rdProc78North),
	.emptyNorth(emptyProc78North),
	.dataInNorth(dataInProc78North),
	.rdSouth(rdProc78South),
	.emptySouth(emptyProc78South),
	.dataInSouth(dataInProc78South),
	.wrSouth(wrProc78South),
	.fullSouth(fullProc78South),
	.dataOutSouth(dataOutProc78South),
	.rdEast(rdProc78East),
	.emptyEast(emptyProc78East),
	.dataInEast(dataInProc78East),
	.wrEast(wrProc78East),
	.fullEast(fullProc78East),
	.dataOutEast(dataOutProc78East));
 
//PROCESSOR 79
system proc79(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe79),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe79),
	.rdNorth(rdProc79North),
	.emptyNorth(emptyProc79North),
	.dataInNorth(dataInProc79North),
	.wrNorth(wrProc79North),
	.fullNorth(fullProc79North),
	.dataOutNorth(dataOutProc79North),
	.rdSouth(rdProc79South),
	.emptySouth(emptyProc79South),
	.dataInSouth(dataInProc79South),
	.wrSouth(wrProc79South),
	.fullSouth(fullProc79South),
	.dataOutSouth(dataOutProc79South),
	.rdEast(rdProc79East),
	.emptyEast(emptyProc79East),
	.dataInEast(dataInProc79East),
	.wrEast(wrProc79East),
	.fullEast(fullProc79East),
	.dataOutEast(dataOutProc79East),
	.rdWest(rdProc79West),
	.emptyWest(emptyProc79West),
	.dataInWest(dataInProc79West),
	.wrWest(wrProc79West),
	.fullWest(fullProc79West),
	.dataOutWest(dataOutProc79West));
 
//PROCESSOR 80
system proc80(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe80),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe80),
	.rdNorth(rdProc80North),
	.emptyNorth(emptyProc80North),
	.dataInNorth(dataInProc80North),
	.wrNorth(wrProc80North),
	.fullNorth(fullProc80North),
	.dataOutNorth(dataOutProc80North),
	.rdSouth(rdProc80South),
	.emptySouth(emptyProc80South),
	.dataInSouth(dataInProc80South),
	.wrSouth(wrProc80South),
	.fullSouth(fullProc80South),
	.dataOutSouth(dataOutProc80South),
	.rdEast(rdProc80East),
	.emptyEast(emptyProc80East),
	.dataInEast(dataInProc80East),
	.wrEast(wrProc80East),
	.fullEast(fullProc80East),
	.dataOutEast(dataOutProc80East),
	.rdWest(rdProc80West),
	.emptyWest(emptyProc80West),
	.dataInWest(dataInProc80West),
	.wrWest(wrProc80West),
	.fullWest(fullProc80West),
	.dataOutWest(dataOutProc80West));
 
//PROCESSOR 81
system proc81(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe81),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe81),
	.rdNorth(rdProc81North),
	.emptyNorth(emptyProc81North),
	.dataInNorth(dataInProc81North),
	.wrNorth(wrProc81North),
	.fullNorth(fullProc81North),
	.dataOutNorth(dataOutProc81North),
	.rdSouth(rdProc81South),
	.emptySouth(emptyProc81South),
	.dataInSouth(dataInProc81South),
	.wrSouth(wrProc81South),
	.fullSouth(fullProc81South),
	.dataOutSouth(dataOutProc81South),
	.rdEast(rdProc81East),
	.emptyEast(emptyProc81East),
	.dataInEast(dataInProc81East),
	.wrEast(wrProc81East),
	.fullEast(fullProc81East),
	.dataOutEast(dataOutProc81East),
	.rdWest(rdProc81West),
	.emptyWest(emptyProc81West),
	.dataInWest(dataInProc81West),
	.wrWest(wrProc81West),
	.fullWest(fullProc81West),
	.dataOutWest(dataOutProc81West));
 
//PROCESSOR 82
system proc82(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe82),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe82),
	.rdNorth(rdProc82North),
	.emptyNorth(emptyProc82North),
	.dataInNorth(dataInProc82North),
	.wrNorth(wrProc82North),
	.fullNorth(fullProc82North),
	.dataOutNorth(dataOutProc82North),
	.rdSouth(rdProc82South),
	.emptySouth(emptyProc82South),
	.dataInSouth(dataInProc82South),
	.wrSouth(wrProc82South),
	.fullSouth(fullProc82South),
	.dataOutSouth(dataOutProc82South),
	.rdEast(rdProc82East),
	.emptyEast(emptyProc82East),
	.dataInEast(dataInProc82East),
	.wrEast(wrProc82East),
	.fullEast(fullProc82East),
	.dataOutEast(dataOutProc82East),
	.rdWest(rdProc82West),
	.emptyWest(emptyProc82West),
	.dataInWest(dataInProc82West),
	.wrWest(wrProc82West),
	.fullWest(fullProc82West),
	.dataOutWest(dataOutProc82West));
 
//PROCESSOR 83
system proc83(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe83),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe83),
	.rdNorth(rdProc83North),
	.emptyNorth(emptyProc83North),
	.dataInNorth(dataInProc83North),
	.wrNorth(wrProc83North),
	.fullNorth(fullProc83North),
	.dataOutNorth(dataOutProc83North),
	.rdSouth(rdProc83South),
	.emptySouth(emptyProc83South),
	.dataInSouth(dataInProc83South),
	.wrSouth(wrProc83South),
	.fullSouth(fullProc83South),
	.dataOutSouth(dataOutProc83South),
	.rdEast(rdProc83East),
	.emptyEast(emptyProc83East),
	.dataInEast(dataInProc83East),
	.wrEast(wrProc83East),
	.fullEast(fullProc83East),
	.dataOutEast(dataOutProc83East),
	.rdWest(rdProc83West),
	.emptyWest(emptyProc83West),
	.dataInWest(dataInProc83West),
	.wrWest(wrProc83West),
	.fullWest(fullProc83West),
	.dataOutWest(dataOutProc83West));
 
//PROCESSOR 84
system proc84(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe84),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe84),
	.rdNorth(rdProc84North),
	.emptyNorth(emptyProc84North),
	.dataInNorth(dataInProc84North),
	.wrNorth(wrProc84North),
	.fullNorth(fullProc84North),
	.dataOutNorth(dataOutProc84North),
	.rdSouth(rdProc84South),
	.emptySouth(emptyProc84South),
	.dataInSouth(dataInProc84South),
	.wrSouth(wrProc84South),
	.fullSouth(fullProc84South),
	.dataOutSouth(dataOutProc84South),
	.rdEast(rdProc84East),
	.emptyEast(emptyProc84East),
	.dataInEast(dataInProc84East),
	.wrEast(wrProc84East),
	.fullEast(fullProc84East),
	.dataOutEast(dataOutProc84East),
	.rdWest(rdProc84West),
	.emptyWest(emptyProc84West),
	.dataInWest(dataInProc84West),
	.wrWest(wrProc84West),
	.fullWest(fullProc84West),
	.dataOutWest(dataOutProc84West));
 
//PROCESSOR 85
system proc85(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe85),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe85),
	.rdNorth(rdProc85North),
	.emptyNorth(emptyProc85North),
	.dataInNorth(dataInProc85North),
	.wrNorth(wrProc85North),
	.fullNorth(fullProc85North),
	.dataOutNorth(dataOutProc85North),
	.rdSouth(rdProc85South),
	.emptySouth(emptyProc85South),
	.dataInSouth(dataInProc85South),
	.wrSouth(wrProc85South),
	.fullSouth(fullProc85South),
	.dataOutSouth(dataOutProc85South),
	.rdEast(rdProc85East),
	.emptyEast(emptyProc85East),
	.dataInEast(dataInProc85East),
	.wrEast(wrProc85East),
	.fullEast(fullProc85East),
	.dataOutEast(dataOutProc85East),
	.rdWest(rdProc85West),
	.emptyWest(emptyProc85West),
	.dataInWest(dataInProc85West),
	.wrWest(wrProc85West),
	.fullWest(fullProc85West),
	.dataOutWest(dataOutProc85West));
 
//PROCESSOR 86
system proc86(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe86),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe86),
	.rdNorth(rdProc86North),
	.emptyNorth(emptyProc86North),
	.dataInNorth(dataInProc86North),
	.wrNorth(wrProc86North),
	.fullNorth(fullProc86North),
	.dataOutNorth(dataOutProc86North),
	.rdSouth(rdProc86South),
	.emptySouth(emptyProc86South),
	.dataInSouth(dataInProc86South),
	.wrSouth(wrProc86South),
	.fullSouth(fullProc86South),
	.dataOutSouth(dataOutProc86South),
	.rdEast(rdProc86East),
	.emptyEast(emptyProc86East),
	.dataInEast(dataInProc86East),
	.wrEast(wrProc86East),
	.fullEast(fullProc86East),
	.dataOutEast(dataOutProc86East),
	.rdWest(rdProc86West),
	.emptyWest(emptyProc86West),
	.dataInWest(dataInProc86West),
	.wrWest(wrProc86West),
	.fullWest(fullProc86West),
	.dataOutWest(dataOutProc86West));
 
//PROCESSOR 87
system proc87(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe87),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe87),
	.rdNorth(rdProc87North),
	.emptyNorth(emptyProc87North),
	.dataInNorth(dataInProc87North),
	.wrNorth(wrProc87North),
	.fullNorth(fullProc87North),
	.dataOutNorth(dataOutProc87North),
	.rdSouth(rdProc87South),
	.emptySouth(emptyProc87South),
	.dataInSouth(dataInProc87South),
	.wrSouth(wrProc87South),
	.fullSouth(fullProc87South),
	.dataOutSouth(dataOutProc87South),
	.rdEast(rdProc87East),
	.emptyEast(emptyProc87East),
	.dataInEast(dataInProc87East),
	.wrEast(wrProc87East),
	.fullEast(fullProc87East),
	.dataOutEast(dataOutProc87East),
	.rdWest(rdProc87West),
	.emptyWest(emptyProc87West),
	.dataInWest(dataInProc87West),
	.wrWest(wrProc87West),
	.fullWest(fullProc87West),
	.dataOutWest(dataOutProc87West));
 
//PROCESSOR 88
system proc88(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe88),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe88),
	.rdNorth(rdProc88North),
	.emptyNorth(emptyProc88North),
	.dataInNorth(dataInProc88North),
	.wrNorth(wrProc88North),
	.fullNorth(fullProc88North),
	.dataOutNorth(dataOutProc88North),
	.rdSouth(rdProc88South),
	.emptySouth(emptyProc88South),
	.dataInSouth(dataInProc88South),
	.wrSouth(wrProc88South),
	.fullSouth(fullProc88South),
	.dataOutSouth(dataOutProc88South),
	.rdEast(rdProc88East),
	.emptyEast(emptyProc88East),
	.dataInEast(dataInProc88East),
	.wrEast(wrProc88East),
	.fullEast(fullProc88East),
	.dataOutEast(dataOutProc88East),
	.rdWest(rdProc88West),
	.emptyWest(emptyProc88West),
	.dataInWest(dataInProc88West),
	.wrWest(wrProc88West),
	.fullWest(fullProc88West),
	.dataOutWest(dataOutProc88West));
 
//PROCESSOR 89
system proc89(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe89),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe89),
	.rdNorth(rdProc89North),
	.emptyNorth(emptyProc89North),
	.dataInNorth(dataInProc89North),
	.wrNorth(wrProc89North),
	.fullNorth(fullProc89North),
	.dataOutNorth(dataOutProc89North),
	.rdSouth(rdProc89South),
	.emptySouth(emptyProc89South),
	.dataInSouth(dataInProc89South),
	.wrSouth(wrProc89South),
	.fullSouth(fullProc89South),
	.dataOutSouth(dataOutProc89South),
	.rdEast(rdProc89East),
	.emptyEast(emptyProc89East),
	.dataInEast(dataInProc89East),
	.wrEast(wrProc89East),
	.fullEast(fullProc89East),
	.dataOutEast(dataOutProc89East),
	.rdWest(rdProc89West),
	.emptyWest(emptyProc89West),
	.dataInWest(dataInProc89West),
	.wrWest(wrProc89West),
	.fullWest(fullProc89West),
	.dataOutWest(dataOutProc89West));
 
//PROCESSOR 90
system proc90(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe90),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe90),
	.rdNorth(rdProc90North),
	.emptyNorth(emptyProc90North),
	.dataInNorth(dataInProc90North),
	.wrNorth(wrProc90North),
	.fullNorth(fullProc90North),
	.dataOutNorth(dataOutProc90North),
	.rdSouth(rdProc90South),
	.emptySouth(emptyProc90South),
	.dataInSouth(dataInProc90South),
	.wrSouth(wrProc90South),
	.fullSouth(fullProc90South),
	.dataOutSouth(dataOutProc90South),
	.rdWest(rdProc90West),
	.emptyWest(emptyProc90West),
	.dataInWest(dataInProc90West),
	.wrWest(wrProc90West),
	.fullWest(fullProc90West),
	.dataOutWest(dataOutProc90West));
 
//PROCESSOR 91
system proc91(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe91),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe91),
	.wrNorth(wrProc91North),
	.fullNorth(fullProc91North),
	.dataOutNorth(dataOutProc91North),
	.rdNorth(rdProc91North),
	.emptyNorth(emptyProc91North),
	.dataInNorth(dataInProc91North),
	.rdSouth(rdProc91South),
	.emptySouth(emptyProc91South),
	.dataInSouth(dataInProc91South),
	.wrSouth(wrProc91South),
	.fullSouth(fullProc91South),
	.dataOutSouth(dataOutProc91South),
	.rdEast(rdProc91East),
	.emptyEast(emptyProc91East),
	.dataInEast(dataInProc91East),
	.wrEast(wrProc91East),
	.fullEast(fullProc91East),
	.dataOutEast(dataOutProc91East));
 
//PROCESSOR 92
system proc92(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe92),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe92),
	.rdNorth(rdProc92North),
	.emptyNorth(emptyProc92North),
	.dataInNorth(dataInProc92North),
	.wrNorth(wrProc92North),
	.fullNorth(fullProc92North),
	.dataOutNorth(dataOutProc92North),
	.rdSouth(rdProc92South),
	.emptySouth(emptyProc92South),
	.dataInSouth(dataInProc92South),
	.wrSouth(wrProc92South),
	.fullSouth(fullProc92South),
	.dataOutSouth(dataOutProc92South),
	.rdEast(rdProc92East),
	.emptyEast(emptyProc92East),
	.dataInEast(dataInProc92East),
	.wrEast(wrProc92East),
	.fullEast(fullProc92East),
	.dataOutEast(dataOutProc92East),
	.rdWest(rdProc92West),
	.emptyWest(emptyProc92West),
	.dataInWest(dataInProc92West),
	.wrWest(wrProc92West),
	.fullWest(fullProc92West),
	.dataOutWest(dataOutProc92West));
 
//PROCESSOR 93
system proc93(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe93),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe93),
	.rdNorth(rdProc93North),
	.emptyNorth(emptyProc93North),
	.dataInNorth(dataInProc93North),
	.wrNorth(wrProc93North),
	.fullNorth(fullProc93North),
	.dataOutNorth(dataOutProc93North),
	.rdSouth(rdProc93South),
	.emptySouth(emptyProc93South),
	.dataInSouth(dataInProc93South),
	.wrSouth(wrProc93South),
	.fullSouth(fullProc93South),
	.dataOutSouth(dataOutProc93South),
	.rdEast(rdProc93East),
	.emptyEast(emptyProc93East),
	.dataInEast(dataInProc93East),
	.wrEast(wrProc93East),
	.fullEast(fullProc93East),
	.dataOutEast(dataOutProc93East),
	.rdWest(rdProc93West),
	.emptyWest(emptyProc93West),
	.dataInWest(dataInProc93West),
	.wrWest(wrProc93West),
	.fullWest(fullProc93West),
	.dataOutWest(dataOutProc93West));
 
//PROCESSOR 94
system proc94(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe94),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe94),
	.rdNorth(rdProc94North),
	.emptyNorth(emptyProc94North),
	.dataInNorth(dataInProc94North),
	.wrNorth(wrProc94North),
	.fullNorth(fullProc94North),
	.dataOutNorth(dataOutProc94North),
	.rdSouth(rdProc94South),
	.emptySouth(emptyProc94South),
	.dataInSouth(dataInProc94South),
	.wrSouth(wrProc94South),
	.fullSouth(fullProc94South),
	.dataOutSouth(dataOutProc94South),
	.rdEast(rdProc94East),
	.emptyEast(emptyProc94East),
	.dataInEast(dataInProc94East),
	.wrEast(wrProc94East),
	.fullEast(fullProc94East),
	.dataOutEast(dataOutProc94East),
	.rdWest(rdProc94West),
	.emptyWest(emptyProc94West),
	.dataInWest(dataInProc94West),
	.wrWest(wrProc94West),
	.fullWest(fullProc94West),
	.dataOutWest(dataOutProc94West));
 
//PROCESSOR 95
system proc95(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe95),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe95),
	.rdNorth(rdProc95North),
	.emptyNorth(emptyProc95North),
	.dataInNorth(dataInProc95North),
	.wrNorth(wrProc95North),
	.fullNorth(fullProc95North),
	.dataOutNorth(dataOutProc95North),
	.rdSouth(rdProc95South),
	.emptySouth(emptyProc95South),
	.dataInSouth(dataInProc95South),
	.wrSouth(wrProc95South),
	.fullSouth(fullProc95South),
	.dataOutSouth(dataOutProc95South),
	.rdEast(rdProc95East),
	.emptyEast(emptyProc95East),
	.dataInEast(dataInProc95East),
	.wrEast(wrProc95East),
	.fullEast(fullProc95East),
	.dataOutEast(dataOutProc95East),
	.rdWest(rdProc95West),
	.emptyWest(emptyProc95West),
	.dataInWest(dataInProc95West),
	.wrWest(wrProc95West),
	.fullWest(fullProc95West),
	.dataOutWest(dataOutProc95West));
 
//PROCESSOR 96
system proc96(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe96),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe96),
	.rdNorth(rdProc96North),
	.emptyNorth(emptyProc96North),
	.dataInNorth(dataInProc96North),
	.wrNorth(wrProc96North),
	.fullNorth(fullProc96North),
	.dataOutNorth(dataOutProc96North),
	.rdSouth(rdProc96South),
	.emptySouth(emptyProc96South),
	.dataInSouth(dataInProc96South),
	.wrSouth(wrProc96South),
	.fullSouth(fullProc96South),
	.dataOutSouth(dataOutProc96South),
	.rdEast(rdProc96East),
	.emptyEast(emptyProc96East),
	.dataInEast(dataInProc96East),
	.wrEast(wrProc96East),
	.fullEast(fullProc96East),
	.dataOutEast(dataOutProc96East),
	.rdWest(rdProc96West),
	.emptyWest(emptyProc96West),
	.dataInWest(dataInProc96West),
	.wrWest(wrProc96West),
	.fullWest(fullProc96West),
	.dataOutWest(dataOutProc96West));
 
//PROCESSOR 97
system proc97(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe97),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe97),
	.rdNorth(rdProc97North),
	.emptyNorth(emptyProc97North),
	.dataInNorth(dataInProc97North),
	.wrNorth(wrProc97North),
	.fullNorth(fullProc97North),
	.dataOutNorth(dataOutProc97North),
	.rdSouth(rdProc97South),
	.emptySouth(emptyProc97South),
	.dataInSouth(dataInProc97South),
	.wrSouth(wrProc97South),
	.fullSouth(fullProc97South),
	.dataOutSouth(dataOutProc97South),
	.rdEast(rdProc97East),
	.emptyEast(emptyProc97East),
	.dataInEast(dataInProc97East),
	.wrEast(wrProc97East),
	.fullEast(fullProc97East),
	.dataOutEast(dataOutProc97East),
	.rdWest(rdProc97West),
	.emptyWest(emptyProc97West),
	.dataInWest(dataInProc97West),
	.wrWest(wrProc97West),
	.fullWest(fullProc97West),
	.dataOutWest(dataOutProc97West));
 
//PROCESSOR 98
system proc98(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe98),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe98),
	.rdNorth(rdProc98North),
	.emptyNorth(emptyProc98North),
	.dataInNorth(dataInProc98North),
	.wrNorth(wrProc98North),
	.fullNorth(fullProc98North),
	.dataOutNorth(dataOutProc98North),
	.rdSouth(rdProc98South),
	.emptySouth(emptyProc98South),
	.dataInSouth(dataInProc98South),
	.wrSouth(wrProc98South),
	.fullSouth(fullProc98South),
	.dataOutSouth(dataOutProc98South),
	.rdEast(rdProc98East),
	.emptyEast(emptyProc98East),
	.dataInEast(dataInProc98East),
	.wrEast(wrProc98East),
	.fullEast(fullProc98East),
	.dataOutEast(dataOutProc98East),
	.rdWest(rdProc98West),
	.emptyWest(emptyProc98West),
	.dataInWest(dataInProc98West),
	.wrWest(wrProc98West),
	.fullWest(fullProc98West),
	.dataOutWest(dataOutProc98West));
 
//PROCESSOR 99
system proc99(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe99),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe99),
	.rdNorth(rdProc99North),
	.emptyNorth(emptyProc99North),
	.dataInNorth(dataInProc99North),
	.wrNorth(wrProc99North),
	.fullNorth(fullProc99North),
	.dataOutNorth(dataOutProc99North),
	.rdSouth(rdProc99South),
	.emptySouth(emptyProc99South),
	.dataInSouth(dataInProc99South),
	.wrSouth(wrProc99South),
	.fullSouth(fullProc99South),
	.dataOutSouth(dataOutProc99South),
	.rdEast(rdProc99East),
	.emptyEast(emptyProc99East),
	.dataInEast(dataInProc99East),
	.wrEast(wrProc99East),
	.fullEast(fullProc99East),
	.dataOutEast(dataOutProc99East),
	.rdWest(rdProc99West),
	.emptyWest(emptyProc99West),
	.dataInWest(dataInProc99West),
	.wrWest(wrProc99West),
	.fullWest(fullProc99West),
	.dataOutWest(dataOutProc99West));
 
//PROCESSOR 100
system proc100(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe100),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe100),
	.rdNorth(rdProc100North),
	.emptyNorth(emptyProc100North),
	.dataInNorth(dataInProc100North),
	.wrNorth(wrProc100North),
	.fullNorth(fullProc100North),
	.dataOutNorth(dataOutProc100North),
	.rdSouth(rdProc100South),
	.emptySouth(emptyProc100South),
	.dataInSouth(dataInProc100South),
	.wrSouth(wrProc100South),
	.fullSouth(fullProc100South),
	.dataOutSouth(dataOutProc100South),
	.rdEast(rdProc100East),
	.emptyEast(emptyProc100East),
	.dataInEast(dataInProc100East),
	.wrEast(wrProc100East),
	.fullEast(fullProc100East),
	.dataOutEast(dataOutProc100East),
	.rdWest(rdProc100West),
	.emptyWest(emptyProc100West),
	.dataInWest(dataInProc100West),
	.wrWest(wrProc100West),
	.fullWest(fullProc100West),
	.dataOutWest(dataOutProc100West));
 
//PROCESSOR 101
system proc101(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe101),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe101),
	.rdNorth(rdProc101North),
	.emptyNorth(emptyProc101North),
	.dataInNorth(dataInProc101North),
	.wrNorth(wrProc101North),
	.fullNorth(fullProc101North),
	.dataOutNorth(dataOutProc101North),
	.rdSouth(rdProc101South),
	.emptySouth(emptyProc101South),
	.dataInSouth(dataInProc101South),
	.wrSouth(wrProc101South),
	.fullSouth(fullProc101South),
	.dataOutSouth(dataOutProc101South),
	.rdEast(rdProc101East),
	.emptyEast(emptyProc101East),
	.dataInEast(dataInProc101East),
	.wrEast(wrProc101East),
	.fullEast(fullProc101East),
	.dataOutEast(dataOutProc101East),
	.rdWest(rdProc101West),
	.emptyWest(emptyProc101West),
	.dataInWest(dataInProc101West),
	.wrWest(wrProc101West),
	.fullWest(fullProc101West),
	.dataOutWest(dataOutProc101West));
 
//PROCESSOR 102
system proc102(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe102),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe102),
	.rdNorth(rdProc102North),
	.emptyNorth(emptyProc102North),
	.dataInNorth(dataInProc102North),
	.wrNorth(wrProc102North),
	.fullNorth(fullProc102North),
	.dataOutNorth(dataOutProc102North),
	.rdSouth(rdProc102South),
	.emptySouth(emptyProc102South),
	.dataInSouth(dataInProc102South),
	.wrSouth(wrProc102South),
	.fullSouth(fullProc102South),
	.dataOutSouth(dataOutProc102South),
	.rdEast(rdProc102East),
	.emptyEast(emptyProc102East),
	.dataInEast(dataInProc102East),
	.wrEast(wrProc102East),
	.fullEast(fullProc102East),
	.dataOutEast(dataOutProc102East),
	.rdWest(rdProc102West),
	.emptyWest(emptyProc102West),
	.dataInWest(dataInProc102West),
	.wrWest(wrProc102West),
	.fullWest(fullProc102West),
	.dataOutWest(dataOutProc102West));
 
//PROCESSOR 103
system proc103(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe103),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe103),
	.rdNorth(rdProc103North),
	.emptyNorth(emptyProc103North),
	.dataInNorth(dataInProc103North),
	.wrNorth(wrProc103North),
	.fullNorth(fullProc103North),
	.dataOutNorth(dataOutProc103North),
	.rdSouth(rdProc103South),
	.emptySouth(emptyProc103South),
	.dataInSouth(dataInProc103South),
	.wrSouth(wrProc103South),
	.fullSouth(fullProc103South),
	.dataOutSouth(dataOutProc103South),
	.rdWest(rdProc103West),
	.emptyWest(emptyProc103West),
	.dataInWest(dataInProc103West),
	.wrWest(wrProc103West),
	.fullWest(fullProc103West),
	.dataOutWest(dataOutProc103West));
 
//PROCESSOR 104
system proc104(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe104),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe104),
	.wrNorth(wrProc104North),
	.fullNorth(fullProc104North),
	.dataOutNorth(dataOutProc104North),
	.rdNorth(rdProc104North),
	.emptyNorth(emptyProc104North),
	.dataInNorth(dataInProc104North),
	.rdSouth(rdProc104South),
	.emptySouth(emptyProc104South),
	.dataInSouth(dataInProc104South),
	.wrSouth(wrProc104South),
	.fullSouth(fullProc104South),
	.dataOutSouth(dataOutProc104South),
	.rdEast(rdProc104East),
	.emptyEast(emptyProc104East),
	.dataInEast(dataInProc104East),
	.wrEast(wrProc104East),
	.fullEast(fullProc104East),
	.dataOutEast(dataOutProc104East));
 
//PROCESSOR 105
system proc105(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe105),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe105),
	.rdNorth(rdProc105North),
	.emptyNorth(emptyProc105North),
	.dataInNorth(dataInProc105North),
	.wrNorth(wrProc105North),
	.fullNorth(fullProc105North),
	.dataOutNorth(dataOutProc105North),
	.rdSouth(rdProc105South),
	.emptySouth(emptyProc105South),
	.dataInSouth(dataInProc105South),
	.wrSouth(wrProc105South),
	.fullSouth(fullProc105South),
	.dataOutSouth(dataOutProc105South),
	.rdEast(rdProc105East),
	.emptyEast(emptyProc105East),
	.dataInEast(dataInProc105East),
	.wrEast(wrProc105East),
	.fullEast(fullProc105East),
	.dataOutEast(dataOutProc105East),
	.rdWest(rdProc105West),
	.emptyWest(emptyProc105West),
	.dataInWest(dataInProc105West),
	.wrWest(wrProc105West),
	.fullWest(fullProc105West),
	.dataOutWest(dataOutProc105West));
 
//PROCESSOR 106
system proc106(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe106),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe106),
	.rdNorth(rdProc106North),
	.emptyNorth(emptyProc106North),
	.dataInNorth(dataInProc106North),
	.wrNorth(wrProc106North),
	.fullNorth(fullProc106North),
	.dataOutNorth(dataOutProc106North),
	.rdSouth(rdProc106South),
	.emptySouth(emptyProc106South),
	.dataInSouth(dataInProc106South),
	.wrSouth(wrProc106South),
	.fullSouth(fullProc106South),
	.dataOutSouth(dataOutProc106South),
	.rdEast(rdProc106East),
	.emptyEast(emptyProc106East),
	.dataInEast(dataInProc106East),
	.wrEast(wrProc106East),
	.fullEast(fullProc106East),
	.dataOutEast(dataOutProc106East),
	.rdWest(rdProc106West),
	.emptyWest(emptyProc106West),
	.dataInWest(dataInProc106West),
	.wrWest(wrProc106West),
	.fullWest(fullProc106West),
	.dataOutWest(dataOutProc106West));
 
//PROCESSOR 107
system proc107(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe107),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe107),
	.rdNorth(rdProc107North),
	.emptyNorth(emptyProc107North),
	.dataInNorth(dataInProc107North),
	.wrNorth(wrProc107North),
	.fullNorth(fullProc107North),
	.dataOutNorth(dataOutProc107North),
	.rdSouth(rdProc107South),
	.emptySouth(emptyProc107South),
	.dataInSouth(dataInProc107South),
	.wrSouth(wrProc107South),
	.fullSouth(fullProc107South),
	.dataOutSouth(dataOutProc107South),
	.rdEast(rdProc107East),
	.emptyEast(emptyProc107East),
	.dataInEast(dataInProc107East),
	.wrEast(wrProc107East),
	.fullEast(fullProc107East),
	.dataOutEast(dataOutProc107East),
	.rdWest(rdProc107West),
	.emptyWest(emptyProc107West),
	.dataInWest(dataInProc107West),
	.wrWest(wrProc107West),
	.fullWest(fullProc107West),
	.dataOutWest(dataOutProc107West));
 
//PROCESSOR 108
system proc108(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe108),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe108),
	.rdNorth(rdProc108North),
	.emptyNorth(emptyProc108North),
	.dataInNorth(dataInProc108North),
	.wrNorth(wrProc108North),
	.fullNorth(fullProc108North),
	.dataOutNorth(dataOutProc108North),
	.rdSouth(rdProc108South),
	.emptySouth(emptyProc108South),
	.dataInSouth(dataInProc108South),
	.wrSouth(wrProc108South),
	.fullSouth(fullProc108South),
	.dataOutSouth(dataOutProc108South),
	.rdEast(rdProc108East),
	.emptyEast(emptyProc108East),
	.dataInEast(dataInProc108East),
	.wrEast(wrProc108East),
	.fullEast(fullProc108East),
	.dataOutEast(dataOutProc108East),
	.rdWest(rdProc108West),
	.emptyWest(emptyProc108West),
	.dataInWest(dataInProc108West),
	.wrWest(wrProc108West),
	.fullWest(fullProc108West),
	.dataOutWest(dataOutProc108West));
 
//PROCESSOR 109
system proc109(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe109),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe109),
	.rdNorth(rdProc109North),
	.emptyNorth(emptyProc109North),
	.dataInNorth(dataInProc109North),
	.wrNorth(wrProc109North),
	.fullNorth(fullProc109North),
	.dataOutNorth(dataOutProc109North),
	.rdSouth(rdProc109South),
	.emptySouth(emptyProc109South),
	.dataInSouth(dataInProc109South),
	.wrSouth(wrProc109South),
	.fullSouth(fullProc109South),
	.dataOutSouth(dataOutProc109South),
	.rdEast(rdProc109East),
	.emptyEast(emptyProc109East),
	.dataInEast(dataInProc109East),
	.wrEast(wrProc109East),
	.fullEast(fullProc109East),
	.dataOutEast(dataOutProc109East),
	.rdWest(rdProc109West),
	.emptyWest(emptyProc109West),
	.dataInWest(dataInProc109West),
	.wrWest(wrProc109West),
	.fullWest(fullProc109West),
	.dataOutWest(dataOutProc109West));
 
//PROCESSOR 110
system proc110(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe110),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe110),
	.rdNorth(rdProc110North),
	.emptyNorth(emptyProc110North),
	.dataInNorth(dataInProc110North),
	.wrNorth(wrProc110North),
	.fullNorth(fullProc110North),
	.dataOutNorth(dataOutProc110North),
	.rdSouth(rdProc110South),
	.emptySouth(emptyProc110South),
	.dataInSouth(dataInProc110South),
	.wrSouth(wrProc110South),
	.fullSouth(fullProc110South),
	.dataOutSouth(dataOutProc110South),
	.rdEast(rdProc110East),
	.emptyEast(emptyProc110East),
	.dataInEast(dataInProc110East),
	.wrEast(wrProc110East),
	.fullEast(fullProc110East),
	.dataOutEast(dataOutProc110East),
	.rdWest(rdProc110West),
	.emptyWest(emptyProc110West),
	.dataInWest(dataInProc110West),
	.wrWest(wrProc110West),
	.fullWest(fullProc110West),
	.dataOutWest(dataOutProc110West));
 
//PROCESSOR 111
system proc111(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe111),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe111),
	.rdNorth(rdProc111North),
	.emptyNorth(emptyProc111North),
	.dataInNorth(dataInProc111North),
	.wrNorth(wrProc111North),
	.fullNorth(fullProc111North),
	.dataOutNorth(dataOutProc111North),
	.rdSouth(rdProc111South),
	.emptySouth(emptyProc111South),
	.dataInSouth(dataInProc111South),
	.wrSouth(wrProc111South),
	.fullSouth(fullProc111South),
	.dataOutSouth(dataOutProc111South),
	.rdEast(rdProc111East),
	.emptyEast(emptyProc111East),
	.dataInEast(dataInProc111East),
	.wrEast(wrProc111East),
	.fullEast(fullProc111East),
	.dataOutEast(dataOutProc111East),
	.rdWest(rdProc111West),
	.emptyWest(emptyProc111West),
	.dataInWest(dataInProc111West),
	.wrWest(wrProc111West),
	.fullWest(fullProc111West),
	.dataOutWest(dataOutProc111West));
 
//PROCESSOR 112
system proc112(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe112),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe112),
	.rdNorth(rdProc112North),
	.emptyNorth(emptyProc112North),
	.dataInNorth(dataInProc112North),
	.wrNorth(wrProc112North),
	.fullNorth(fullProc112North),
	.dataOutNorth(dataOutProc112North),
	.rdSouth(rdProc112South),
	.emptySouth(emptyProc112South),
	.dataInSouth(dataInProc112South),
	.wrSouth(wrProc112South),
	.fullSouth(fullProc112South),
	.dataOutSouth(dataOutProc112South),
	.rdEast(rdProc112East),
	.emptyEast(emptyProc112East),
	.dataInEast(dataInProc112East),
	.wrEast(wrProc112East),
	.fullEast(fullProc112East),
	.dataOutEast(dataOutProc112East),
	.rdWest(rdProc112West),
	.emptyWest(emptyProc112West),
	.dataInWest(dataInProc112West),
	.wrWest(wrProc112West),
	.fullWest(fullProc112West),
	.dataOutWest(dataOutProc112West));
 
//PROCESSOR 113
system proc113(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe113),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe113),
	.rdNorth(rdProc113North),
	.emptyNorth(emptyProc113North),
	.dataInNorth(dataInProc113North),
	.wrNorth(wrProc113North),
	.fullNorth(fullProc113North),
	.dataOutNorth(dataOutProc113North),
	.rdSouth(rdProc113South),
	.emptySouth(emptyProc113South),
	.dataInSouth(dataInProc113South),
	.wrSouth(wrProc113South),
	.fullSouth(fullProc113South),
	.dataOutSouth(dataOutProc113South),
	.rdEast(rdProc113East),
	.emptyEast(emptyProc113East),
	.dataInEast(dataInProc113East),
	.wrEast(wrProc113East),
	.fullEast(fullProc113East),
	.dataOutEast(dataOutProc113East),
	.rdWest(rdProc113West),
	.emptyWest(emptyProc113West),
	.dataInWest(dataInProc113West),
	.wrWest(wrProc113West),
	.fullWest(fullProc113West),
	.dataOutWest(dataOutProc113West));
 
//PROCESSOR 114
system proc114(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe114),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe114),
	.rdNorth(rdProc114North),
	.emptyNorth(emptyProc114North),
	.dataInNorth(dataInProc114North),
	.wrNorth(wrProc114North),
	.fullNorth(fullProc114North),
	.dataOutNorth(dataOutProc114North),
	.rdSouth(rdProc114South),
	.emptySouth(emptyProc114South),
	.dataInSouth(dataInProc114South),
	.wrSouth(wrProc114South),
	.fullSouth(fullProc114South),
	.dataOutSouth(dataOutProc114South),
	.rdEast(rdProc114East),
	.emptyEast(emptyProc114East),
	.dataInEast(dataInProc114East),
	.wrEast(wrProc114East),
	.fullEast(fullProc114East),
	.dataOutEast(dataOutProc114East),
	.rdWest(rdProc114West),
	.emptyWest(emptyProc114West),
	.dataInWest(dataInProc114West),
	.wrWest(wrProc114West),
	.fullWest(fullProc114West),
	.dataOutWest(dataOutProc114West));
 
//PROCESSOR 115
system proc115(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe115),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe115),
	.rdNorth(rdProc115North),
	.emptyNorth(emptyProc115North),
	.dataInNorth(dataInProc115North),
	.wrNorth(wrProc115North),
	.fullNorth(fullProc115North),
	.dataOutNorth(dataOutProc115North),
	.rdSouth(rdProc115South),
	.emptySouth(emptyProc115South),
	.dataInSouth(dataInProc115South),
	.wrSouth(wrProc115South),
	.fullSouth(fullProc115South),
	.dataOutSouth(dataOutProc115South),
	.rdEast(rdProc115East),
	.emptyEast(emptyProc115East),
	.dataInEast(dataInProc115East),
	.wrEast(wrProc115East),
	.fullEast(fullProc115East),
	.dataOutEast(dataOutProc115East),
	.rdWest(rdProc115West),
	.emptyWest(emptyProc115West),
	.dataInWest(dataInProc115West),
	.wrWest(wrProc115West),
	.fullWest(fullProc115West),
	.dataOutWest(dataOutProc115West));
 
//PROCESSOR 116
system proc116(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe116),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe116),
	.rdNorth(rdProc116North),
	.emptyNorth(emptyProc116North),
	.dataInNorth(dataInProc116North),
	.wrNorth(wrProc116North),
	.fullNorth(fullProc116North),
	.dataOutNorth(dataOutProc116North),
	.rdSouth(rdProc116South),
	.emptySouth(emptyProc116South),
	.dataInSouth(dataInProc116South),
	.wrSouth(wrProc116South),
	.fullSouth(fullProc116South),
	.dataOutSouth(dataOutProc116South),
	.rdWest(rdProc116West),
	.emptyWest(emptyProc116West),
	.dataInWest(dataInProc116West),
	.wrWest(wrProc116West),
	.fullWest(fullProc116West),
	.dataOutWest(dataOutProc116West));
 
//PROCESSOR 117
system proc117(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe117),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe117),
	.wrNorth(wrProc117North),
	.fullNorth(fullProc117North),
	.dataOutNorth(dataOutProc117North),
	.rdNorth(rdProc117North),
	.emptyNorth(emptyProc117North),
	.dataInNorth(dataInProc117North),
	.rdSouth(rdProc117South),
	.emptySouth(emptyProc117South),
	.dataInSouth(dataInProc117South),
	.wrSouth(wrProc117South),
	.fullSouth(fullProc117South),
	.dataOutSouth(dataOutProc117South),
	.rdEast(rdProc117East),
	.emptyEast(emptyProc117East),
	.dataInEast(dataInProc117East),
	.wrEast(wrProc117East),
	.fullEast(fullProc117East),
	.dataOutEast(dataOutProc117East));
 
//PROCESSOR 118
system proc118(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe118),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe118),
	.rdNorth(rdProc118North),
	.emptyNorth(emptyProc118North),
	.dataInNorth(dataInProc118North),
	.wrNorth(wrProc118North),
	.fullNorth(fullProc118North),
	.dataOutNorth(dataOutProc118North),
	.rdSouth(rdProc118South),
	.emptySouth(emptyProc118South),
	.dataInSouth(dataInProc118South),
	.wrSouth(wrProc118South),
	.fullSouth(fullProc118South),
	.dataOutSouth(dataOutProc118South),
	.rdEast(rdProc118East),
	.emptyEast(emptyProc118East),
	.dataInEast(dataInProc118East),
	.wrEast(wrProc118East),
	.fullEast(fullProc118East),
	.dataOutEast(dataOutProc118East),
	.rdWest(rdProc118West),
	.emptyWest(emptyProc118West),
	.dataInWest(dataInProc118West),
	.wrWest(wrProc118West),
	.fullWest(fullProc118West),
	.dataOutWest(dataOutProc118West));
 
//PROCESSOR 119
system proc119(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe119),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe119),
	.rdNorth(rdProc119North),
	.emptyNorth(emptyProc119North),
	.dataInNorth(dataInProc119North),
	.wrNorth(wrProc119North),
	.fullNorth(fullProc119North),
	.dataOutNorth(dataOutProc119North),
	.rdSouth(rdProc119South),
	.emptySouth(emptyProc119South),
	.dataInSouth(dataInProc119South),
	.wrSouth(wrProc119South),
	.fullSouth(fullProc119South),
	.dataOutSouth(dataOutProc119South),
	.rdEast(rdProc119East),
	.emptyEast(emptyProc119East),
	.dataInEast(dataInProc119East),
	.wrEast(wrProc119East),
	.fullEast(fullProc119East),
	.dataOutEast(dataOutProc119East),
	.rdWest(rdProc119West),
	.emptyWest(emptyProc119West),
	.dataInWest(dataInProc119West),
	.wrWest(wrProc119West),
	.fullWest(fullProc119West),
	.dataOutWest(dataOutProc119West));
 
//PROCESSOR 120
system proc120(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe120),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe120),
	.rdNorth(rdProc120North),
	.emptyNorth(emptyProc120North),
	.dataInNorth(dataInProc120North),
	.wrNorth(wrProc120North),
	.fullNorth(fullProc120North),
	.dataOutNorth(dataOutProc120North),
	.rdSouth(rdProc120South),
	.emptySouth(emptyProc120South),
	.dataInSouth(dataInProc120South),
	.wrSouth(wrProc120South),
	.fullSouth(fullProc120South),
	.dataOutSouth(dataOutProc120South),
	.rdEast(rdProc120East),
	.emptyEast(emptyProc120East),
	.dataInEast(dataInProc120East),
	.wrEast(wrProc120East),
	.fullEast(fullProc120East),
	.dataOutEast(dataOutProc120East),
	.rdWest(rdProc120West),
	.emptyWest(emptyProc120West),
	.dataInWest(dataInProc120West),
	.wrWest(wrProc120West),
	.fullWest(fullProc120West),
	.dataOutWest(dataOutProc120West));
 
//PROCESSOR 121
system proc121(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe121),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe121),
	.rdNorth(rdProc121North),
	.emptyNorth(emptyProc121North),
	.dataInNorth(dataInProc121North),
	.wrNorth(wrProc121North),
	.fullNorth(fullProc121North),
	.dataOutNorth(dataOutProc121North),
	.rdSouth(rdProc121South),
	.emptySouth(emptyProc121South),
	.dataInSouth(dataInProc121South),
	.wrSouth(wrProc121South),
	.fullSouth(fullProc121South),
	.dataOutSouth(dataOutProc121South),
	.rdEast(rdProc121East),
	.emptyEast(emptyProc121East),
	.dataInEast(dataInProc121East),
	.wrEast(wrProc121East),
	.fullEast(fullProc121East),
	.dataOutEast(dataOutProc121East),
	.rdWest(rdProc121West),
	.emptyWest(emptyProc121West),
	.dataInWest(dataInProc121West),
	.wrWest(wrProc121West),
	.fullWest(fullProc121West),
	.dataOutWest(dataOutProc121West));
 
//PROCESSOR 122
system proc122(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe122),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe122),
	.rdNorth(rdProc122North),
	.emptyNorth(emptyProc122North),
	.dataInNorth(dataInProc122North),
	.wrNorth(wrProc122North),
	.fullNorth(fullProc122North),
	.dataOutNorth(dataOutProc122North),
	.rdSouth(rdProc122South),
	.emptySouth(emptyProc122South),
	.dataInSouth(dataInProc122South),
	.wrSouth(wrProc122South),
	.fullSouth(fullProc122South),
	.dataOutSouth(dataOutProc122South),
	.rdEast(rdProc122East),
	.emptyEast(emptyProc122East),
	.dataInEast(dataInProc122East),
	.wrEast(wrProc122East),
	.fullEast(fullProc122East),
	.dataOutEast(dataOutProc122East),
	.rdWest(rdProc122West),
	.emptyWest(emptyProc122West),
	.dataInWest(dataInProc122West),
	.wrWest(wrProc122West),
	.fullWest(fullProc122West),
	.dataOutWest(dataOutProc122West));
 
//PROCESSOR 123
system proc123(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe123),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe123),
	.rdNorth(rdProc123North),
	.emptyNorth(emptyProc123North),
	.dataInNorth(dataInProc123North),
	.wrNorth(wrProc123North),
	.fullNorth(fullProc123North),
	.dataOutNorth(dataOutProc123North),
	.rdSouth(rdProc123South),
	.emptySouth(emptyProc123South),
	.dataInSouth(dataInProc123South),
	.wrSouth(wrProc123South),
	.fullSouth(fullProc123South),
	.dataOutSouth(dataOutProc123South),
	.rdEast(rdProc123East),
	.emptyEast(emptyProc123East),
	.dataInEast(dataInProc123East),
	.wrEast(wrProc123East),
	.fullEast(fullProc123East),
	.dataOutEast(dataOutProc123East),
	.rdWest(rdProc123West),
	.emptyWest(emptyProc123West),
	.dataInWest(dataInProc123West),
	.wrWest(wrProc123West),
	.fullWest(fullProc123West),
	.dataOutWest(dataOutProc123West));
 
//PROCESSOR 124
system proc124(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe124),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe124),
	.rdNorth(rdProc124North),
	.emptyNorth(emptyProc124North),
	.dataInNorth(dataInProc124North),
	.wrNorth(wrProc124North),
	.fullNorth(fullProc124North),
	.dataOutNorth(dataOutProc124North),
	.rdSouth(rdProc124South),
	.emptySouth(emptyProc124South),
	.dataInSouth(dataInProc124South),
	.wrSouth(wrProc124South),
	.fullSouth(fullProc124South),
	.dataOutSouth(dataOutProc124South),
	.rdEast(rdProc124East),
	.emptyEast(emptyProc124East),
	.dataInEast(dataInProc124East),
	.wrEast(wrProc124East),
	.fullEast(fullProc124East),
	.dataOutEast(dataOutProc124East),
	.rdWest(rdProc124West),
	.emptyWest(emptyProc124West),
	.dataInWest(dataInProc124West),
	.wrWest(wrProc124West),
	.fullWest(fullProc124West),
	.dataOutWest(dataOutProc124West));
 
//PROCESSOR 125
system proc125(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe125),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe125),
	.rdNorth(rdProc125North),
	.emptyNorth(emptyProc125North),
	.dataInNorth(dataInProc125North),
	.wrNorth(wrProc125North),
	.fullNorth(fullProc125North),
	.dataOutNorth(dataOutProc125North),
	.rdSouth(rdProc125South),
	.emptySouth(emptyProc125South),
	.dataInSouth(dataInProc125South),
	.wrSouth(wrProc125South),
	.fullSouth(fullProc125South),
	.dataOutSouth(dataOutProc125South),
	.rdEast(rdProc125East),
	.emptyEast(emptyProc125East),
	.dataInEast(dataInProc125East),
	.wrEast(wrProc125East),
	.fullEast(fullProc125East),
	.dataOutEast(dataOutProc125East),
	.rdWest(rdProc125West),
	.emptyWest(emptyProc125West),
	.dataInWest(dataInProc125West),
	.wrWest(wrProc125West),
	.fullWest(fullProc125West),
	.dataOutWest(dataOutProc125West));
 
//PROCESSOR 126
system proc126(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe126),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe126),
	.rdNorth(rdProc126North),
	.emptyNorth(emptyProc126North),
	.dataInNorth(dataInProc126North),
	.wrNorth(wrProc126North),
	.fullNorth(fullProc126North),
	.dataOutNorth(dataOutProc126North),
	.rdSouth(rdProc126South),
	.emptySouth(emptyProc126South),
	.dataInSouth(dataInProc126South),
	.wrSouth(wrProc126South),
	.fullSouth(fullProc126South),
	.dataOutSouth(dataOutProc126South),
	.rdEast(rdProc126East),
	.emptyEast(emptyProc126East),
	.dataInEast(dataInProc126East),
	.wrEast(wrProc126East),
	.fullEast(fullProc126East),
	.dataOutEast(dataOutProc126East),
	.rdWest(rdProc126West),
	.emptyWest(emptyProc126West),
	.dataInWest(dataInProc126West),
	.wrWest(wrProc126West),
	.fullWest(fullProc126West),
	.dataOutWest(dataOutProc126West));
 
//PROCESSOR 127
system proc127(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe127),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe127),
	.rdNorth(rdProc127North),
	.emptyNorth(emptyProc127North),
	.dataInNorth(dataInProc127North),
	.wrNorth(wrProc127North),
	.fullNorth(fullProc127North),
	.dataOutNorth(dataOutProc127North),
	.rdSouth(rdProc127South),
	.emptySouth(emptyProc127South),
	.dataInSouth(dataInProc127South),
	.wrSouth(wrProc127South),
	.fullSouth(fullProc127South),
	.dataOutSouth(dataOutProc127South),
	.rdEast(rdProc127East),
	.emptyEast(emptyProc127East),
	.dataInEast(dataInProc127East),
	.wrEast(wrProc127East),
	.fullEast(fullProc127East),
	.dataOutEast(dataOutProc127East),
	.rdWest(rdProc127West),
	.emptyWest(emptyProc127West),
	.dataInWest(dataInProc127West),
	.wrWest(wrProc127West),
	.fullWest(fullProc127West),
	.dataOutWest(dataOutProc127West));
 
//PROCESSOR 128
system proc128(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe128),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe128),
	.rdNorth(rdProc128North),
	.emptyNorth(emptyProc128North),
	.dataInNorth(dataInProc128North),
	.wrNorth(wrProc128North),
	.fullNorth(fullProc128North),
	.dataOutNorth(dataOutProc128North),
	.rdSouth(rdProc128South),
	.emptySouth(emptyProc128South),
	.dataInSouth(dataInProc128South),
	.wrSouth(wrProc128South),
	.fullSouth(fullProc128South),
	.dataOutSouth(dataOutProc128South),
	.rdEast(rdProc128East),
	.emptyEast(emptyProc128East),
	.dataInEast(dataInProc128East),
	.wrEast(wrProc128East),
	.fullEast(fullProc128East),
	.dataOutEast(dataOutProc128East),
	.rdWest(rdProc128West),
	.emptyWest(emptyProc128West),
	.dataInWest(dataInProc128West),
	.wrWest(wrProc128West),
	.fullWest(fullProc128West),
	.dataOutWest(dataOutProc128West));
 
//PROCESSOR 129
system proc129(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe129),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe129),
	.rdNorth(rdProc129North),
	.emptyNorth(emptyProc129North),
	.dataInNorth(dataInProc129North),
	.wrNorth(wrProc129North),
	.fullNorth(fullProc129North),
	.dataOutNorth(dataOutProc129North),
	.rdSouth(rdProc129South),
	.emptySouth(emptyProc129South),
	.dataInSouth(dataInProc129South),
	.wrSouth(wrProc129South),
	.fullSouth(fullProc129South),
	.dataOutSouth(dataOutProc129South),
	.rdWest(rdProc129West),
	.emptyWest(emptyProc129West),
	.dataInWest(dataInProc129West),
	.wrWest(wrProc129West),
	.fullWest(fullProc129West),
	.dataOutWest(dataOutProc129West));
 
//PROCESSOR 130
system proc130(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe130),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe130),
	.wrNorth(wrProc130North),
	.fullNorth(fullProc130North),
	.dataOutNorth(dataOutProc130North),
	.rdNorth(rdProc130North),
	.emptyNorth(emptyProc130North),
	.dataInNorth(dataInProc130North),
	.rdSouth(rdProc130South),
	.emptySouth(emptyProc130South),
	.dataInSouth(dataInProc130South),
	.wrSouth(wrProc130South),
	.fullSouth(fullProc130South),
	.dataOutSouth(dataOutProc130South),
	.rdEast(rdProc130East),
	.emptyEast(emptyProc130East),
	.dataInEast(dataInProc130East),
	.wrEast(wrProc130East),
	.fullEast(fullProc130East),
	.dataOutEast(dataOutProc130East));
 
//PROCESSOR 131
system proc131(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe131),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe131),
	.rdNorth(rdProc131North),
	.emptyNorth(emptyProc131North),
	.dataInNorth(dataInProc131North),
	.wrNorth(wrProc131North),
	.fullNorth(fullProc131North),
	.dataOutNorth(dataOutProc131North),
	.rdSouth(rdProc131South),
	.emptySouth(emptyProc131South),
	.dataInSouth(dataInProc131South),
	.wrSouth(wrProc131South),
	.fullSouth(fullProc131South),
	.dataOutSouth(dataOutProc131South),
	.rdEast(rdProc131East),
	.emptyEast(emptyProc131East),
	.dataInEast(dataInProc131East),
	.wrEast(wrProc131East),
	.fullEast(fullProc131East),
	.dataOutEast(dataOutProc131East),
	.rdWest(rdProc131West),
	.emptyWest(emptyProc131West),
	.dataInWest(dataInProc131West),
	.wrWest(wrProc131West),
	.fullWest(fullProc131West),
	.dataOutWest(dataOutProc131West));
 
//PROCESSOR 132
system proc132(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe132),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe132),
	.rdNorth(rdProc132North),
	.emptyNorth(emptyProc132North),
	.dataInNorth(dataInProc132North),
	.wrNorth(wrProc132North),
	.fullNorth(fullProc132North),
	.dataOutNorth(dataOutProc132North),
	.rdSouth(rdProc132South),
	.emptySouth(emptyProc132South),
	.dataInSouth(dataInProc132South),
	.wrSouth(wrProc132South),
	.fullSouth(fullProc132South),
	.dataOutSouth(dataOutProc132South),
	.rdEast(rdProc132East),
	.emptyEast(emptyProc132East),
	.dataInEast(dataInProc132East),
	.wrEast(wrProc132East),
	.fullEast(fullProc132East),
	.dataOutEast(dataOutProc132East),
	.rdWest(rdProc132West),
	.emptyWest(emptyProc132West),
	.dataInWest(dataInProc132West),
	.wrWest(wrProc132West),
	.fullWest(fullProc132West),
	.dataOutWest(dataOutProc132West));
 
//PROCESSOR 133
system proc133(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe133),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe133),
	.rdNorth(rdProc133North),
	.emptyNorth(emptyProc133North),
	.dataInNorth(dataInProc133North),
	.wrNorth(wrProc133North),
	.fullNorth(fullProc133North),
	.dataOutNorth(dataOutProc133North),
	.rdSouth(rdProc133South),
	.emptySouth(emptyProc133South),
	.dataInSouth(dataInProc133South),
	.wrSouth(wrProc133South),
	.fullSouth(fullProc133South),
	.dataOutSouth(dataOutProc133South),
	.rdEast(rdProc133East),
	.emptyEast(emptyProc133East),
	.dataInEast(dataInProc133East),
	.wrEast(wrProc133East),
	.fullEast(fullProc133East),
	.dataOutEast(dataOutProc133East),
	.rdWest(rdProc133West),
	.emptyWest(emptyProc133West),
	.dataInWest(dataInProc133West),
	.wrWest(wrProc133West),
	.fullWest(fullProc133West),
	.dataOutWest(dataOutProc133West));
 
//PROCESSOR 134
system proc134(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe134),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe134),
	.rdNorth(rdProc134North),
	.emptyNorth(emptyProc134North),
	.dataInNorth(dataInProc134North),
	.wrNorth(wrProc134North),
	.fullNorth(fullProc134North),
	.dataOutNorth(dataOutProc134North),
	.rdSouth(rdProc134South),
	.emptySouth(emptyProc134South),
	.dataInSouth(dataInProc134South),
	.wrSouth(wrProc134South),
	.fullSouth(fullProc134South),
	.dataOutSouth(dataOutProc134South),
	.rdEast(rdProc134East),
	.emptyEast(emptyProc134East),
	.dataInEast(dataInProc134East),
	.wrEast(wrProc134East),
	.fullEast(fullProc134East),
	.dataOutEast(dataOutProc134East),
	.rdWest(rdProc134West),
	.emptyWest(emptyProc134West),
	.dataInWest(dataInProc134West),
	.wrWest(wrProc134West),
	.fullWest(fullProc134West),
	.dataOutWest(dataOutProc134West));
 
//PROCESSOR 135
system proc135(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe135),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe135),
	.rdNorth(rdProc135North),
	.emptyNorth(emptyProc135North),
	.dataInNorth(dataInProc135North),
	.wrNorth(wrProc135North),
	.fullNorth(fullProc135North),
	.dataOutNorth(dataOutProc135North),
	.rdSouth(rdProc135South),
	.emptySouth(emptyProc135South),
	.dataInSouth(dataInProc135South),
	.wrSouth(wrProc135South),
	.fullSouth(fullProc135South),
	.dataOutSouth(dataOutProc135South),
	.rdEast(rdProc135East),
	.emptyEast(emptyProc135East),
	.dataInEast(dataInProc135East),
	.wrEast(wrProc135East),
	.fullEast(fullProc135East),
	.dataOutEast(dataOutProc135East),
	.rdWest(rdProc135West),
	.emptyWest(emptyProc135West),
	.dataInWest(dataInProc135West),
	.wrWest(wrProc135West),
	.fullWest(fullProc135West),
	.dataOutWest(dataOutProc135West));
 
//PROCESSOR 136
system proc136(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe136),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe136),
	.rdNorth(rdProc136North),
	.emptyNorth(emptyProc136North),
	.dataInNorth(dataInProc136North),
	.wrNorth(wrProc136North),
	.fullNorth(fullProc136North),
	.dataOutNorth(dataOutProc136North),
	.rdSouth(rdProc136South),
	.emptySouth(emptyProc136South),
	.dataInSouth(dataInProc136South),
	.wrSouth(wrProc136South),
	.fullSouth(fullProc136South),
	.dataOutSouth(dataOutProc136South),
	.rdEast(rdProc136East),
	.emptyEast(emptyProc136East),
	.dataInEast(dataInProc136East),
	.wrEast(wrProc136East),
	.fullEast(fullProc136East),
	.dataOutEast(dataOutProc136East),
	.rdWest(rdProc136West),
	.emptyWest(emptyProc136West),
	.dataInWest(dataInProc136West),
	.wrWest(wrProc136West),
	.fullWest(fullProc136West),
	.dataOutWest(dataOutProc136West));
 
//PROCESSOR 137
system proc137(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe137),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe137),
	.rdNorth(rdProc137North),
	.emptyNorth(emptyProc137North),
	.dataInNorth(dataInProc137North),
	.wrNorth(wrProc137North),
	.fullNorth(fullProc137North),
	.dataOutNorth(dataOutProc137North),
	.rdSouth(rdProc137South),
	.emptySouth(emptyProc137South),
	.dataInSouth(dataInProc137South),
	.wrSouth(wrProc137South),
	.fullSouth(fullProc137South),
	.dataOutSouth(dataOutProc137South),
	.rdEast(rdProc137East),
	.emptyEast(emptyProc137East),
	.dataInEast(dataInProc137East),
	.wrEast(wrProc137East),
	.fullEast(fullProc137East),
	.dataOutEast(dataOutProc137East),
	.rdWest(rdProc137West),
	.emptyWest(emptyProc137West),
	.dataInWest(dataInProc137West),
	.wrWest(wrProc137West),
	.fullWest(fullProc137West),
	.dataOutWest(dataOutProc137West));
 
//PROCESSOR 138
system proc138(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe138),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe138),
	.rdNorth(rdProc138North),
	.emptyNorth(emptyProc138North),
	.dataInNorth(dataInProc138North),
	.wrNorth(wrProc138North),
	.fullNorth(fullProc138North),
	.dataOutNorth(dataOutProc138North),
	.rdSouth(rdProc138South),
	.emptySouth(emptyProc138South),
	.dataInSouth(dataInProc138South),
	.wrSouth(wrProc138South),
	.fullSouth(fullProc138South),
	.dataOutSouth(dataOutProc138South),
	.rdEast(rdProc138East),
	.emptyEast(emptyProc138East),
	.dataInEast(dataInProc138East),
	.wrEast(wrProc138East),
	.fullEast(fullProc138East),
	.dataOutEast(dataOutProc138East),
	.rdWest(rdProc138West),
	.emptyWest(emptyProc138West),
	.dataInWest(dataInProc138West),
	.wrWest(wrProc138West),
	.fullWest(fullProc138West),
	.dataOutWest(dataOutProc138West));
 
//PROCESSOR 139
system proc139(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe139),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe139),
	.rdNorth(rdProc139North),
	.emptyNorth(emptyProc139North),
	.dataInNorth(dataInProc139North),
	.wrNorth(wrProc139North),
	.fullNorth(fullProc139North),
	.dataOutNorth(dataOutProc139North),
	.rdSouth(rdProc139South),
	.emptySouth(emptyProc139South),
	.dataInSouth(dataInProc139South),
	.wrSouth(wrProc139South),
	.fullSouth(fullProc139South),
	.dataOutSouth(dataOutProc139South),
	.rdEast(rdProc139East),
	.emptyEast(emptyProc139East),
	.dataInEast(dataInProc139East),
	.wrEast(wrProc139East),
	.fullEast(fullProc139East),
	.dataOutEast(dataOutProc139East),
	.rdWest(rdProc139West),
	.emptyWest(emptyProc139West),
	.dataInWest(dataInProc139West),
	.wrWest(wrProc139West),
	.fullWest(fullProc139West),
	.dataOutWest(dataOutProc139West));
 
//PROCESSOR 140
system proc140(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe140),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe140),
	.rdNorth(rdProc140North),
	.emptyNorth(emptyProc140North),
	.dataInNorth(dataInProc140North),
	.wrNorth(wrProc140North),
	.fullNorth(fullProc140North),
	.dataOutNorth(dataOutProc140North),
	.rdSouth(rdProc140South),
	.emptySouth(emptyProc140South),
	.dataInSouth(dataInProc140South),
	.wrSouth(wrProc140South),
	.fullSouth(fullProc140South),
	.dataOutSouth(dataOutProc140South),
	.rdEast(rdProc140East),
	.emptyEast(emptyProc140East),
	.dataInEast(dataInProc140East),
	.wrEast(wrProc140East),
	.fullEast(fullProc140East),
	.dataOutEast(dataOutProc140East),
	.rdWest(rdProc140West),
	.emptyWest(emptyProc140West),
	.dataInWest(dataInProc140West),
	.wrWest(wrProc140West),
	.fullWest(fullProc140West),
	.dataOutWest(dataOutProc140West));
 
//PROCESSOR 141
system proc141(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe141),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe141),
	.rdNorth(rdProc141North),
	.emptyNorth(emptyProc141North),
	.dataInNorth(dataInProc141North),
	.wrNorth(wrProc141North),
	.fullNorth(fullProc141North),
	.dataOutNorth(dataOutProc141North),
	.rdSouth(rdProc141South),
	.emptySouth(emptyProc141South),
	.dataInSouth(dataInProc141South),
	.wrSouth(wrProc141South),
	.fullSouth(fullProc141South),
	.dataOutSouth(dataOutProc141South),
	.rdEast(rdProc141East),
	.emptyEast(emptyProc141East),
	.dataInEast(dataInProc141East),
	.wrEast(wrProc141East),
	.fullEast(fullProc141East),
	.dataOutEast(dataOutProc141East),
	.rdWest(rdProc141West),
	.emptyWest(emptyProc141West),
	.dataInWest(dataInProc141West),
	.wrWest(wrProc141West),
	.fullWest(fullProc141West),
	.dataOutWest(dataOutProc141West));
 
//PROCESSOR 142
system proc142(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe142),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe142),
	.rdNorth(rdProc142North),
	.emptyNorth(emptyProc142North),
	.dataInNorth(dataInProc142North),
	.wrNorth(wrProc142North),
	.fullNorth(fullProc142North),
	.dataOutNorth(dataOutProc142North),
	.rdSouth(rdProc142South),
	.emptySouth(emptyProc142South),
	.dataInSouth(dataInProc142South),
	.wrSouth(wrProc142South),
	.fullSouth(fullProc142South),
	.dataOutSouth(dataOutProc142South),
	.rdWest(rdProc142West),
	.emptyWest(emptyProc142West),
	.dataInWest(dataInProc142West),
	.wrWest(wrProc142West),
	.fullWest(fullProc142West),
	.dataOutWest(dataOutProc142West));
 
//PROCESSOR 143
system proc143(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe143),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe143),
	.rdNorth(rdProc143North),
	.emptyNorth(emptyProc143North),
	.dataInNorth(dataInProc143North),
	.wrNorth(wrProc143North),
	.fullNorth(fullProc143North),
	.dataOutNorth(dataOutProc143North),
	.rdEast(rdProc143East),
	.emptyEast(emptyProc143East),
	.dataInEast(dataInProc143East),
	.wrEast(wrProc143East),
	.fullEast(fullProc143East),
	.dataOutEast(dataOutProc143East));
 
//PROCESSOR 144
system proc144(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe144),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe144),
	.rdNorth(rdProc144North),
	.emptyNorth(emptyProc144North),
	.dataInNorth(dataInProc144North),
	.wrNorth(wrProc144North),
	.fullNorth(fullProc144North),
	.dataOutNorth(dataOutProc144North),
	.rdEast(rdProc144East),
	.emptyEast(emptyProc144East),
	.dataInEast(dataInProc144East),
	.wrEast(wrProc144East),
	.fullEast(fullProc144East),
	.dataOutEast(dataOutProc144East),
	.rdWest(rdProc144West),
	.emptyWest(emptyProc144West),
	.dataInWest(dataInProc144West),
	.wrWest(wrProc144West),
	.fullWest(fullProc144West),
	.dataOutWest(dataOutProc144West));
 
//PROCESSOR 145
system proc145(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe145),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe145),
	.rdNorth(rdProc145North),
	.emptyNorth(emptyProc145North),
	.dataInNorth(dataInProc145North),
	.wrNorth(wrProc145North),
	.fullNorth(fullProc145North),
	.dataOutNorth(dataOutProc145North),
	.rdEast(rdProc145East),
	.emptyEast(emptyProc145East),
	.dataInEast(dataInProc145East),
	.wrEast(wrProc145East),
	.fullEast(fullProc145East),
	.dataOutEast(dataOutProc145East),
	.rdWest(rdProc145West),
	.emptyWest(emptyProc145West),
	.dataInWest(dataInProc145West),
	.wrWest(wrProc145West),
	.fullWest(fullProc145West),
	.dataOutWest(dataOutProc145West));
 
//PROCESSOR 146
system proc146(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe146),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe146),
	.rdNorth(rdProc146North),
	.emptyNorth(emptyProc146North),
	.dataInNorth(dataInProc146North),
	.wrNorth(wrProc146North),
	.fullNorth(fullProc146North),
	.dataOutNorth(dataOutProc146North),
	.rdEast(rdProc146East),
	.emptyEast(emptyProc146East),
	.dataInEast(dataInProc146East),
	.wrEast(wrProc146East),
	.fullEast(fullProc146East),
	.dataOutEast(dataOutProc146East),
	.rdWest(rdProc146West),
	.emptyWest(emptyProc146West),
	.dataInWest(dataInProc146West),
	.wrWest(wrProc146West),
	.fullWest(fullProc146West),
	.dataOutWest(dataOutProc146West));
 
//PROCESSOR 147
system proc147(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe147),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe147),
	.rdNorth(rdProc147North),
	.emptyNorth(emptyProc147North),
	.dataInNorth(dataInProc147North),
	.wrNorth(wrProc147North),
	.fullNorth(fullProc147North),
	.dataOutNorth(dataOutProc147North),
	.rdEast(rdProc147East),
	.emptyEast(emptyProc147East),
	.dataInEast(dataInProc147East),
	.wrEast(wrProc147East),
	.fullEast(fullProc147East),
	.dataOutEast(dataOutProc147East),
	.rdWest(rdProc147West),
	.emptyWest(emptyProc147West),
	.dataInWest(dataInProc147West),
	.wrWest(wrProc147West),
	.fullWest(fullProc147West),
	.dataOutWest(dataOutProc147West));
 
//PROCESSOR 148
system proc148(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe148),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe148),
	.rdNorth(rdProc148North),
	.emptyNorth(emptyProc148North),
	.dataInNorth(dataInProc148North),
	.wrNorth(wrProc148North),
	.fullNorth(fullProc148North),
	.dataOutNorth(dataOutProc148North),
	.rdEast(rdProc148East),
	.emptyEast(emptyProc148East),
	.dataInEast(dataInProc148East),
	.wrEast(wrProc148East),
	.fullEast(fullProc148East),
	.dataOutEast(dataOutProc148East),
	.rdWest(rdProc148West),
	.emptyWest(emptyProc148West),
	.dataInWest(dataInProc148West),
	.wrWest(wrProc148West),
	.fullWest(fullProc148West),
	.dataOutWest(dataOutProc148West));
 
//PROCESSOR 149
system proc149(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe149),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe149),
	.rdNorth(rdProc149North),
	.emptyNorth(emptyProc149North),
	.dataInNorth(dataInProc149North),
	.wrNorth(wrProc149North),
	.fullNorth(fullProc149North),
	.dataOutNorth(dataOutProc149North),
	.rdEast(rdProc149East),
	.emptyEast(emptyProc149East),
	.dataInEast(dataInProc149East),
	.wrEast(wrProc149East),
	.fullEast(fullProc149East),
	.dataOutEast(dataOutProc149East),
	.rdWest(rdProc149West),
	.emptyWest(emptyProc149West),
	.dataInWest(dataInProc149West),
	.wrWest(wrProc149West),
	.fullWest(fullProc149West),
	.dataOutWest(dataOutProc149West));
 
//PROCESSOR 150
system proc150(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe150),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe150),
	.rdNorth(rdProc150North),
	.emptyNorth(emptyProc150North),
	.dataInNorth(dataInProc150North),
	.wrNorth(wrProc150North),
	.fullNorth(fullProc150North),
	.dataOutNorth(dataOutProc150North),
	.rdEast(rdProc150East),
	.emptyEast(emptyProc150East),
	.dataInEast(dataInProc150East),
	.wrEast(wrProc150East),
	.fullEast(fullProc150East),
	.dataOutEast(dataOutProc150East),
	.rdWest(rdProc150West),
	.emptyWest(emptyProc150West),
	.dataInWest(dataInProc150West),
	.wrWest(wrProc150West),
	.fullWest(fullProc150West),
	.dataOutWest(dataOutProc150West));
 
//PROCESSOR 151
system proc151(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe151),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe151),
	.rdNorth(rdProc151North),
	.emptyNorth(emptyProc151North),
	.dataInNorth(dataInProc151North),
	.wrNorth(wrProc151North),
	.fullNorth(fullProc151North),
	.dataOutNorth(dataOutProc151North),
	.rdEast(rdProc151East),
	.emptyEast(emptyProc151East),
	.dataInEast(dataInProc151East),
	.wrEast(wrProc151East),
	.fullEast(fullProc151East),
	.dataOutEast(dataOutProc151East),
	.rdWest(rdProc151West),
	.emptyWest(emptyProc151West),
	.dataInWest(dataInProc151West),
	.wrWest(wrProc151West),
	.fullWest(fullProc151West),
	.dataOutWest(dataOutProc151West));
 
//PROCESSOR 152
system proc152(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe152),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe152),
	.rdNorth(rdProc152North),
	.emptyNorth(emptyProc152North),
	.dataInNorth(dataInProc152North),
	.wrNorth(wrProc152North),
	.fullNorth(fullProc152North),
	.dataOutNorth(dataOutProc152North),
	.rdEast(rdProc152East),
	.emptyEast(emptyProc152East),
	.dataInEast(dataInProc152East),
	.wrEast(wrProc152East),
	.fullEast(fullProc152East),
	.dataOutEast(dataOutProc152East),
	.rdWest(rdProc152West),
	.emptyWest(emptyProc152West),
	.dataInWest(dataInProc152West),
	.wrWest(wrProc152West),
	.fullWest(fullProc152West),
	.dataOutWest(dataOutProc152West));
 
//PROCESSOR 153
system proc153(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe153),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe153),
	.rdNorth(rdProc153North),
	.emptyNorth(emptyProc153North),
	.dataInNorth(dataInProc153North),
	.wrNorth(wrProc153North),
	.fullNorth(fullProc153North),
	.dataOutNorth(dataOutProc153North),
	.rdEast(rdProc153East),
	.emptyEast(emptyProc153East),
	.dataInEast(dataInProc153East),
	.wrEast(wrProc153East),
	.fullEast(fullProc153East),
	.dataOutEast(dataOutProc153East),
	.rdWest(rdProc153West),
	.emptyWest(emptyProc153West),
	.dataInWest(dataInProc153West),
	.wrWest(wrProc153West),
	.fullWest(fullProc153West),
	.dataOutWest(dataOutProc153West));
 
//PROCESSOR 154
system proc154(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe154),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe154),
	.rdNorth(rdProc154North),
	.emptyNorth(emptyProc154North),
	.dataInNorth(dataInProc154North),
	.wrNorth(wrProc154North),
	.fullNorth(fullProc154North),
	.dataOutNorth(dataOutProc154North),
	.rdEast(rdProc154East),
	.emptyEast(emptyProc154East),
	.dataInEast(dataInProc154East),
	.wrEast(wrProc154East),
	.fullEast(fullProc154East),
	.dataOutEast(dataOutProc154East),
	.rdWest(rdProc154West),
	.emptyWest(emptyProc154West),
	.dataInWest(dataInProc154West),
	.wrWest(wrProc154West),
	.fullWest(fullProc154West),
	.dataOutWest(dataOutProc154West));
 
//PROCESSOR 155
system proc155(.clk(clk),
	.resetn (resetn),
	.boot_iaddr(boot_iaddr),
	.boot_idata(boot_idata),
	.boot_iwe(boot_iwe155),
	.boot_daddr(boot_daddr),
	.boot_ddata(boot_ddata),
	.boot_dwe(boot_dwe155),
	.rdNorth(rdProc155North),
	.emptyNorth(emptyProc155North),
	.dataInNorth(dataInProc155North),
	.wrNorth(wrProc155North),
	.fullNorth(fullProc155North),
	.dataOutNorth(dataOutProc155North),
	.wrWest(wrProc155West),
	.fullWest(fullProc155West),
	.dataOutWest(dataOutProc155West),
	.rdWest(rdProc155West),
	.emptyWest(emptyProc155West),
	.dataInWest(dataInProc155West));
	
	//FIFO 1 TO 0 
fifo fifo_proc1_to_proc0(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc1West),
	.full(fullProc1West),
	.dataIn(dataOutProc1West),
	.rd(rdProc0East),
	.empty(emptyProc0East),
	.dataOut(dataInProc0East));
	
	//FIFO 0 TO 1
fifo fifo_proc0_to_proc1(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc0East),
	.full(fullProc0East),
	.dataIn(dataOutProc0East),
	.rd(rdProc1West),
	.empty(emptyProc1West),
	.dataOut(dataInProc1West));
	
	//FIFO 2 TO 1 
fifo fifo_proc2_to_proc1(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc2West),
	.full(fullProc2West),
	.dataIn(dataOutProc2West),
	.rd(rdProc1East),
	.empty(emptyProc1East),
	.dataOut(dataInProc1East));
	
	//FIFO 1 TO 2
fifo fifo_proc1_to_proc2(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc1East),
	.full(fullProc1East),
	.dataIn(dataOutProc1East),
	.rd(rdProc2West),
	.empty(emptyProc2West),
	.dataOut(dataInProc2West));
	
	//FIFO 3 TO 2 
fifo fifo_proc3_to_proc2(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc3West),
	.full(fullProc3West),
	.dataIn(dataOutProc3West),
	.rd(rdProc2East),
	.empty(emptyProc2East),
	.dataOut(dataInProc2East));
	
	//FIFO 2 TO 3
fifo fifo_proc2_to_proc3(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc2East),
	.full(fullProc2East),
	.dataIn(dataOutProc2East),
	.rd(rdProc3West),
	.empty(emptyProc3West),
	.dataOut(dataInProc3West));
	
	//FIFO 4 TO 3 
fifo fifo_proc4_to_proc3(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc4West),
	.full(fullProc4West),
	.dataIn(dataOutProc4West),
	.rd(rdProc3East),
	.empty(emptyProc3East),
	.dataOut(dataInProc3East));
	
	//FIFO 3 TO 4
fifo fifo_proc3_to_proc4(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc3East),
	.full(fullProc3East),
	.dataIn(dataOutProc3East),
	.rd(rdProc4West),
	.empty(emptyProc4West),
	.dataOut(dataInProc4West));
	
	//FIFO 5 TO 4 
fifo fifo_proc5_to_proc4(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc5West),
	.full(fullProc5West),
	.dataIn(dataOutProc5West),
	.rd(rdProc4East),
	.empty(emptyProc4East),
	.dataOut(dataInProc4East));
	
	//FIFO 4 TO 5
fifo fifo_proc4_to_proc5(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc4East),
	.full(fullProc4East),
	.dataIn(dataOutProc4East),
	.rd(rdProc5West),
	.empty(emptyProc5West),
	.dataOut(dataInProc5West));
	
	//FIFO 6 TO 5 
fifo fifo_proc6_to_proc5(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc6West),
	.full(fullProc6West),
	.dataIn(dataOutProc6West),
	.rd(rdProc5East),
	.empty(emptyProc5East),
	.dataOut(dataInProc5East));
	
	//FIFO 5 TO 6
fifo fifo_proc5_to_proc6(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc5East),
	.full(fullProc5East),
	.dataIn(dataOutProc5East),
	.rd(rdProc6West),
	.empty(emptyProc6West),
	.dataOut(dataInProc6West));
	
	//FIFO 7 TO 6 
fifo fifo_proc7_to_proc6(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc7West),
	.full(fullProc7West),
	.dataIn(dataOutProc7West),
	.rd(rdProc6East),
	.empty(emptyProc6East),
	.dataOut(dataInProc6East));
	
	//FIFO 6 TO 7
fifo fifo_proc6_to_proc7(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc6East),
	.full(fullProc6East),
	.dataIn(dataOutProc6East),
	.rd(rdProc7West),
	.empty(emptyProc7West),
	.dataOut(dataInProc7West));
	
	//FIFO 8 TO 7 
fifo fifo_proc8_to_proc7(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc8West),
	.full(fullProc8West),
	.dataIn(dataOutProc8West),
	.rd(rdProc7East),
	.empty(emptyProc7East),
	.dataOut(dataInProc7East));
	
	//FIFO 7 TO 8
fifo fifo_proc7_to_proc8(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc7East),
	.full(fullProc7East),
	.dataIn(dataOutProc7East),
	.rd(rdProc8West),
	.empty(emptyProc8West),
	.dataOut(dataInProc8West));
	
	//FIFO 9 TO 8 
fifo fifo_proc9_to_proc8(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc9West),
	.full(fullProc9West),
	.dataIn(dataOutProc9West),
	.rd(rdProc8East),
	.empty(emptyProc8East),
	.dataOut(dataInProc8East));
	
	//FIFO 8 TO 9
fifo fifo_proc8_to_proc9(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc8East),
	.full(fullProc8East),
	.dataIn(dataOutProc8East),
	.rd(rdProc9West),
	.empty(emptyProc9West),
	.dataOut(dataInProc9West));
	
	//FIFO 10 TO 9 
fifo fifo_proc10_to_proc9(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc10West),
	.full(fullProc10West),
	.dataIn(dataOutProc10West),
	.rd(rdProc9East),
	.empty(emptyProc9East),
	.dataOut(dataInProc9East));
	
	//FIFO 9 TO 10
fifo fifo_proc9_to_proc10(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc9East),
	.full(fullProc9East),
	.dataIn(dataOutProc9East),
	.rd(rdProc10West),
	.empty(emptyProc10West),
	.dataOut(dataInProc10West));
	
	//FIFO 11 TO 10 
fifo fifo_proc11_to_proc10(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc11West),
	.full(fullProc11West),
	.dataIn(dataOutProc11West),
	.rd(rdProc10East),
	.empty(emptyProc10East),
	.dataOut(dataInProc10East));
	
	//FIFO 10 TO 11
fifo fifo_proc10_to_proc11(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc10East),
	.full(fullProc10East),
	.dataIn(dataOutProc10East),
	.rd(rdProc11West),
	.empty(emptyProc11West),
	.dataOut(dataInProc11West));
	
	//FIFO 12 TO 11 
fifo fifo_proc12_to_proc11(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc12West),
	.full(fullProc12West),
	.dataIn(dataOutProc12West),
	.rd(rdProc11East),
	.empty(emptyProc11East),
	.dataOut(dataInProc11East));
	
	//FIFO 11 TO 12
fifo fifo_proc11_to_proc12(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc11East),
	.full(fullProc11East),
	.dataIn(dataOutProc11East),
	.rd(rdProc12West),
	.empty(emptyProc12West),
	.dataOut(dataInProc12West));

	//FIFO 13 TO 0 
fifo fifo_proc13_to_proc0(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc13North),
	.full(fullProc13North),
	.dataIn(dataOutProc13North),
	.rd(rdProc0South),
	.empty(emptyProc0South),
	.dataOut(dataInProc0South));
	
	//FIFO 0 TO 13
fifo fifo_proc0_to_proc13(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc0South),
	.full(fullProc0South),
	.dataIn(dataOutProc0South),
	.rd(rdProc13North),
	.empty(emptyProc13North),
	.dataOut(dataInProc13North));

	//FIFO 14 TO 13 
fifo fifo_proc14_to_proc13(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc14West),
	.full(fullProc14West),
	.dataIn(dataOutProc14West),
	.rd(rdProc13East),
	.empty(emptyProc13East),
	.dataOut(dataInProc13East));
	
	//FIFO 13 TO 14
fifo fifo_proc13_to_proc14(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc13East),
	.full(fullProc13East),
	.dataIn(dataOutProc13East),
	.rd(rdProc14West),
	.empty(emptyProc14West),
	.dataOut(dataInProc14West));
	
	//FIFO 14 TO 1 
fifo fifo_proc14_to_proc1(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc14North),
	.full(fullProc14North),
	.dataIn(dataOutProc14North),
	.rd(rdProc1South),
	.empty(emptyProc1South),
	.dataOut(dataInProc1South));
	
	//FIFO 1 TO 14
fifo fifo_proc1_to_proc14(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc1South),
	.full(fullProc1South),
	.dataIn(dataOutProc1South),
	.rd(rdProc14North),
	.empty(emptyProc14North),
	.dataOut(dataInProc14North));

	//FIFO 15 TO 14 
fifo fifo_proc15_to_proc14(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc15West),
	.full(fullProc15West),
	.dataIn(dataOutProc15West),
	.rd(rdProc14East),
	.empty(emptyProc14East),
	.dataOut(dataInProc14East));
	
	//FIFO 14 TO 15
fifo fifo_proc14_to_proc15(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc14East),
	.full(fullProc14East),
	.dataIn(dataOutProc14East),
	.rd(rdProc15West),
	.empty(emptyProc15West),
	.dataOut(dataInProc15West));
	
	//FIFO 15 TO 2 
fifo fifo_proc15_to_proc2(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc15North),
	.full(fullProc15North),
	.dataIn(dataOutProc15North),
	.rd(rdProc2South),
	.empty(emptyProc2South),
	.dataOut(dataInProc2South));
	
	//FIFO 2 TO 15
fifo fifo_proc2_to_proc15(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc2South),
	.full(fullProc2South),
	.dataIn(dataOutProc2South),
	.rd(rdProc15North),
	.empty(emptyProc15North),
	.dataOut(dataInProc15North));

	//FIFO 16 TO 15 
fifo fifo_proc16_to_proc15(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc16West),
	.full(fullProc16West),
	.dataIn(dataOutProc16West),
	.rd(rdProc15East),
	.empty(emptyProc15East),
	.dataOut(dataInProc15East));
	
	//FIFO 15 TO 16
fifo fifo_proc15_to_proc16(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc15East),
	.full(fullProc15East),
	.dataIn(dataOutProc15East),
	.rd(rdProc16West),
	.empty(emptyProc16West),
	.dataOut(dataInProc16West));
	
	//FIFO 16 TO 3 
fifo fifo_proc16_to_proc3(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc16North),
	.full(fullProc16North),
	.dataIn(dataOutProc16North),
	.rd(rdProc3South),
	.empty(emptyProc3South),
	.dataOut(dataInProc3South));
	
	//FIFO 3 TO 16
fifo fifo_proc3_to_proc16(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc3South),
	.full(fullProc3South),
	.dataIn(dataOutProc3South),
	.rd(rdProc16North),
	.empty(emptyProc16North),
	.dataOut(dataInProc16North));

	//FIFO 17 TO 16 
fifo fifo_proc17_to_proc16(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc17West),
	.full(fullProc17West),
	.dataIn(dataOutProc17West),
	.rd(rdProc16East),
	.empty(emptyProc16East),
	.dataOut(dataInProc16East));
	
	//FIFO 16 TO 17
fifo fifo_proc16_to_proc17(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc16East),
	.full(fullProc16East),
	.dataIn(dataOutProc16East),
	.rd(rdProc17West),
	.empty(emptyProc17West),
	.dataOut(dataInProc17West));
	
	//FIFO 17 TO 4 
fifo fifo_proc17_to_proc4(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc17North),
	.full(fullProc17North),
	.dataIn(dataOutProc17North),
	.rd(rdProc4South),
	.empty(emptyProc4South),
	.dataOut(dataInProc4South));
	
	//FIFO 4 TO 17
fifo fifo_proc4_to_proc17(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc4South),
	.full(fullProc4South),
	.dataIn(dataOutProc4South),
	.rd(rdProc17North),
	.empty(emptyProc17North),
	.dataOut(dataInProc17North));

	//FIFO 18 TO 17 
fifo fifo_proc18_to_proc17(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc18West),
	.full(fullProc18West),
	.dataIn(dataOutProc18West),
	.rd(rdProc17East),
	.empty(emptyProc17East),
	.dataOut(dataInProc17East));
	
	//FIFO 17 TO 18
fifo fifo_proc17_to_proc18(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc17East),
	.full(fullProc17East),
	.dataIn(dataOutProc17East),
	.rd(rdProc18West),
	.empty(emptyProc18West),
	.dataOut(dataInProc18West));
	
	//FIFO 18 TO 5 
fifo fifo_proc18_to_proc5(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc18North),
	.full(fullProc18North),
	.dataIn(dataOutProc18North),
	.rd(rdProc5South),
	.empty(emptyProc5South),
	.dataOut(dataInProc5South));
	
	//FIFO 5 TO 18
fifo fifo_proc5_to_proc18(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc5South),
	.full(fullProc5South),
	.dataIn(dataOutProc5South),
	.rd(rdProc18North),
	.empty(emptyProc18North),
	.dataOut(dataInProc18North));

	//FIFO 19 TO 18 
fifo fifo_proc19_to_proc18(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc19West),
	.full(fullProc19West),
	.dataIn(dataOutProc19West),
	.rd(rdProc18East),
	.empty(emptyProc18East),
	.dataOut(dataInProc18East));
	
	//FIFO 18 TO 19
fifo fifo_proc18_to_proc19(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc18East),
	.full(fullProc18East),
	.dataIn(dataOutProc18East),
	.rd(rdProc19West),
	.empty(emptyProc19West),
	.dataOut(dataInProc19West));
	
	//FIFO 19 TO 6 
fifo fifo_proc19_to_proc6(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc19North),
	.full(fullProc19North),
	.dataIn(dataOutProc19North),
	.rd(rdProc6South),
	.empty(emptyProc6South),
	.dataOut(dataInProc6South));
	
	//FIFO 6 TO 19
fifo fifo_proc6_to_proc19(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc6South),
	.full(fullProc6South),
	.dataIn(dataOutProc6South),
	.rd(rdProc19North),
	.empty(emptyProc19North),
	.dataOut(dataInProc19North));

	//FIFO 20 TO 19 
fifo fifo_proc20_to_proc19(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc20West),
	.full(fullProc20West),
	.dataIn(dataOutProc20West),
	.rd(rdProc19East),
	.empty(emptyProc19East),
	.dataOut(dataInProc19East));
	
	//FIFO 19 TO 20
fifo fifo_proc19_to_proc20(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc19East),
	.full(fullProc19East),
	.dataIn(dataOutProc19East),
	.rd(rdProc20West),
	.empty(emptyProc20West),
	.dataOut(dataInProc20West));
	
	//FIFO 20 TO 7 
fifo fifo_proc20_to_proc7(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc20North),
	.full(fullProc20North),
	.dataIn(dataOutProc20North),
	.rd(rdProc7South),
	.empty(emptyProc7South),
	.dataOut(dataInProc7South));
	
	//FIFO 7 TO 20
fifo fifo_proc7_to_proc20(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc7South),
	.full(fullProc7South),
	.dataIn(dataOutProc7South),
	.rd(rdProc20North),
	.empty(emptyProc20North),
	.dataOut(dataInProc20North));

	//FIFO 21 TO 20 
fifo fifo_proc21_to_proc20(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc21West),
	.full(fullProc21West),
	.dataIn(dataOutProc21West),
	.rd(rdProc20East),
	.empty(emptyProc20East),
	.dataOut(dataInProc20East));
	
	//FIFO 20 TO 21
fifo fifo_proc20_to_proc21(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc20East),
	.full(fullProc20East),
	.dataIn(dataOutProc20East),
	.rd(rdProc21West),
	.empty(emptyProc21West),
	.dataOut(dataInProc21West));
	
	//FIFO 21 TO 8 
fifo fifo_proc21_to_proc8(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc21North),
	.full(fullProc21North),
	.dataIn(dataOutProc21North),
	.rd(rdProc8South),
	.empty(emptyProc8South),
	.dataOut(dataInProc8South));
	
	//FIFO 8 TO 21
fifo fifo_proc8_to_proc21(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc8South),
	.full(fullProc8South),
	.dataIn(dataOutProc8South),
	.rd(rdProc21North),
	.empty(emptyProc21North),
	.dataOut(dataInProc21North));

	//FIFO 22 TO 21 
fifo fifo_proc22_to_proc21(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc22West),
	.full(fullProc22West),
	.dataIn(dataOutProc22West),
	.rd(rdProc21East),
	.empty(emptyProc21East),
	.dataOut(dataInProc21East));
	
	//FIFO 21 TO 22
fifo fifo_proc21_to_proc22(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc21East),
	.full(fullProc21East),
	.dataIn(dataOutProc21East),
	.rd(rdProc22West),
	.empty(emptyProc22West),
	.dataOut(dataInProc22West));
	
	//FIFO 22 TO 9 
fifo fifo_proc22_to_proc9(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc22North),
	.full(fullProc22North),
	.dataIn(dataOutProc22North),
	.rd(rdProc9South),
	.empty(emptyProc9South),
	.dataOut(dataInProc9South));
	
	//FIFO 9 TO 22
fifo fifo_proc9_to_proc22(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc9South),
	.full(fullProc9South),
	.dataIn(dataOutProc9South),
	.rd(rdProc22North),
	.empty(emptyProc22North),
	.dataOut(dataInProc22North));

	//FIFO 23 TO 22 
fifo fifo_proc23_to_proc22(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc23West),
	.full(fullProc23West),
	.dataIn(dataOutProc23West),
	.rd(rdProc22East),
	.empty(emptyProc22East),
	.dataOut(dataInProc22East));
	
	//FIFO 22 TO 23
fifo fifo_proc22_to_proc23(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc22East),
	.full(fullProc22East),
	.dataIn(dataOutProc22East),
	.rd(rdProc23West),
	.empty(emptyProc23West),
	.dataOut(dataInProc23West));
	
	//FIFO 23 TO 10 
fifo fifo_proc23_to_proc10(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc23North),
	.full(fullProc23North),
	.dataIn(dataOutProc23North),
	.rd(rdProc10South),
	.empty(emptyProc10South),
	.dataOut(dataInProc10South));
	
	//FIFO 10 TO 23
fifo fifo_proc10_to_proc23(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc10South),
	.full(fullProc10South),
	.dataIn(dataOutProc10South),
	.rd(rdProc23North),
	.empty(emptyProc23North),
	.dataOut(dataInProc23North));

	//FIFO 24 TO 23 
fifo fifo_proc24_to_proc23(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc24West),
	.full(fullProc24West),
	.dataIn(dataOutProc24West),
	.rd(rdProc23East),
	.empty(emptyProc23East),
	.dataOut(dataInProc23East));
	
	//FIFO 23 TO 24
fifo fifo_proc23_to_proc24(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc23East),
	.full(fullProc23East),
	.dataIn(dataOutProc23East),
	.rd(rdProc24West),
	.empty(emptyProc24West),
	.dataOut(dataInProc24West));
	
	//FIFO 24 TO 11 
fifo fifo_proc24_to_proc11(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc24North),
	.full(fullProc24North),
	.dataIn(dataOutProc24North),
	.rd(rdProc11South),
	.empty(emptyProc11South),
	.dataOut(dataInProc11South));
	
	//FIFO 11 TO 24
fifo fifo_proc11_to_proc24(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc11South),
	.full(fullProc11South),
	.dataIn(dataOutProc11South),
	.rd(rdProc24North),
	.empty(emptyProc24North),
	.dataOut(dataInProc24North));

	//FIFO 25 TO 24 
fifo fifo_proc25_to_proc24(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc25West),
	.full(fullProc25West),
	.dataIn(dataOutProc25West),
	.rd(rdProc24East),
	.empty(emptyProc24East),
	.dataOut(dataInProc24East));
	
	//FIFO 24 TO 25
fifo fifo_proc24_to_proc25(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc24East),
	.full(fullProc24East),
	.dataIn(dataOutProc24East),
	.rd(rdProc25West),
	.empty(emptyProc25West),
	.dataOut(dataInProc25West));
	
	//FIFO 25 TO 12 
fifo fifo_proc25_to_proc12(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc25North),
	.full(fullProc25North),
	.dataIn(dataOutProc25North),
	.rd(rdProc12South),
	.empty(emptyProc12South),
	.dataOut(dataInProc12South));
	
	//FIFO 12 TO 25
fifo fifo_proc12_to_proc25(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc12South),
	.full(fullProc12South),
	.dataIn(dataOutProc12South),
	.rd(rdProc25North),
	.empty(emptyProc25North),
	.dataOut(dataInProc25North));

	//FIFO 26 TO 13 
fifo fifo_proc26_to_proc13(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc26North),
	.full(fullProc26North),
	.dataIn(dataOutProc26North),
	.rd(rdProc13South),
	.empty(emptyProc13South),
	.dataOut(dataInProc13South));
	
	//FIFO 13 TO 26
fifo fifo_proc13_to_proc26(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc13South),
	.full(fullProc13South),
	.dataIn(dataOutProc13South),
	.rd(rdProc26North),
	.empty(emptyProc26North),
	.dataOut(dataInProc26North));

	//FIFO 27 TO 26 
fifo fifo_proc27_to_proc26(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc27West),
	.full(fullProc27West),
	.dataIn(dataOutProc27West),
	.rd(rdProc26East),
	.empty(emptyProc26East),
	.dataOut(dataInProc26East));
	
	//FIFO 26 TO 27
fifo fifo_proc26_to_proc27(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc26East),
	.full(fullProc26East),
	.dataIn(dataOutProc26East),
	.rd(rdProc27West),
	.empty(emptyProc27West),
	.dataOut(dataInProc27West));
	
	//FIFO 27 TO 14 
fifo fifo_proc27_to_proc14(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc27North),
	.full(fullProc27North),
	.dataIn(dataOutProc27North),
	.rd(rdProc14South),
	.empty(emptyProc14South),
	.dataOut(dataInProc14South));
	
	//FIFO 14 TO 27
fifo fifo_proc14_to_proc27(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc14South),
	.full(fullProc14South),
	.dataIn(dataOutProc14South),
	.rd(rdProc27North),
	.empty(emptyProc27North),
	.dataOut(dataInProc27North));

	//FIFO 28 TO 27 
fifo fifo_proc28_to_proc27(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc28West),
	.full(fullProc28West),
	.dataIn(dataOutProc28West),
	.rd(rdProc27East),
	.empty(emptyProc27East),
	.dataOut(dataInProc27East));
	
	//FIFO 27 TO 28
fifo fifo_proc27_to_proc28(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc27East),
	.full(fullProc27East),
	.dataIn(dataOutProc27East),
	.rd(rdProc28West),
	.empty(emptyProc28West),
	.dataOut(dataInProc28West));
	
	//FIFO 28 TO 15 
fifo fifo_proc28_to_proc15(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc28North),
	.full(fullProc28North),
	.dataIn(dataOutProc28North),
	.rd(rdProc15South),
	.empty(emptyProc15South),
	.dataOut(dataInProc15South));
	
	//FIFO 15 TO 28
fifo fifo_proc15_to_proc28(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc15South),
	.full(fullProc15South),
	.dataIn(dataOutProc15South),
	.rd(rdProc28North),
	.empty(emptyProc28North),
	.dataOut(dataInProc28North));

	//FIFO 29 TO 28 
fifo fifo_proc29_to_proc28(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc29West),
	.full(fullProc29West),
	.dataIn(dataOutProc29West),
	.rd(rdProc28East),
	.empty(emptyProc28East),
	.dataOut(dataInProc28East));
	
	//FIFO 28 TO 29
fifo fifo_proc28_to_proc29(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc28East),
	.full(fullProc28East),
	.dataIn(dataOutProc28East),
	.rd(rdProc29West),
	.empty(emptyProc29West),
	.dataOut(dataInProc29West));
	
	//FIFO 29 TO 16 
fifo fifo_proc29_to_proc16(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc29North),
	.full(fullProc29North),
	.dataIn(dataOutProc29North),
	.rd(rdProc16South),
	.empty(emptyProc16South),
	.dataOut(dataInProc16South));
	
	//FIFO 16 TO 29
fifo fifo_proc16_to_proc29(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc16South),
	.full(fullProc16South),
	.dataIn(dataOutProc16South),
	.rd(rdProc29North),
	.empty(emptyProc29North),
	.dataOut(dataInProc29North));

	//FIFO 30 TO 29 
fifo fifo_proc30_to_proc29(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc30West),
	.full(fullProc30West),
	.dataIn(dataOutProc30West),
	.rd(rdProc29East),
	.empty(emptyProc29East),
	.dataOut(dataInProc29East));
	
	//FIFO 29 TO 30
fifo fifo_proc29_to_proc30(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc29East),
	.full(fullProc29East),
	.dataIn(dataOutProc29East),
	.rd(rdProc30West),
	.empty(emptyProc30West),
	.dataOut(dataInProc30West));
	
	//FIFO 30 TO 17 
fifo fifo_proc30_to_proc17(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc30North),
	.full(fullProc30North),
	.dataIn(dataOutProc30North),
	.rd(rdProc17South),
	.empty(emptyProc17South),
	.dataOut(dataInProc17South));
	
	//FIFO 17 TO 30
fifo fifo_proc17_to_proc30(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc17South),
	.full(fullProc17South),
	.dataIn(dataOutProc17South),
	.rd(rdProc30North),
	.empty(emptyProc30North),
	.dataOut(dataInProc30North));

	//FIFO 31 TO 30 
fifo fifo_proc31_to_proc30(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc31West),
	.full(fullProc31West),
	.dataIn(dataOutProc31West),
	.rd(rdProc30East),
	.empty(emptyProc30East),
	.dataOut(dataInProc30East));
	
	//FIFO 30 TO 31
fifo fifo_proc30_to_proc31(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc30East),
	.full(fullProc30East),
	.dataIn(dataOutProc30East),
	.rd(rdProc31West),
	.empty(emptyProc31West),
	.dataOut(dataInProc31West));
	
	//FIFO 31 TO 18 
fifo fifo_proc31_to_proc18(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc31North),
	.full(fullProc31North),
	.dataIn(dataOutProc31North),
	.rd(rdProc18South),
	.empty(emptyProc18South),
	.dataOut(dataInProc18South));
	
	//FIFO 18 TO 31
fifo fifo_proc18_to_proc31(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc18South),
	.full(fullProc18South),
	.dataIn(dataOutProc18South),
	.rd(rdProc31North),
	.empty(emptyProc31North),
	.dataOut(dataInProc31North));

	//FIFO 32 TO 31 
fifo fifo_proc32_to_proc31(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc32West),
	.full(fullProc32West),
	.dataIn(dataOutProc32West),
	.rd(rdProc31East),
	.empty(emptyProc31East),
	.dataOut(dataInProc31East));
	
	//FIFO 31 TO 32
fifo fifo_proc31_to_proc32(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc31East),
	.full(fullProc31East),
	.dataIn(dataOutProc31East),
	.rd(rdProc32West),
	.empty(emptyProc32West),
	.dataOut(dataInProc32West));
	
	//FIFO 32 TO 19 
fifo fifo_proc32_to_proc19(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc32North),
	.full(fullProc32North),
	.dataIn(dataOutProc32North),
	.rd(rdProc19South),
	.empty(emptyProc19South),
	.dataOut(dataInProc19South));
	
	//FIFO 19 TO 32
fifo fifo_proc19_to_proc32(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc19South),
	.full(fullProc19South),
	.dataIn(dataOutProc19South),
	.rd(rdProc32North),
	.empty(emptyProc32North),
	.dataOut(dataInProc32North));

	//FIFO 33 TO 32 
fifo fifo_proc33_to_proc32(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc33West),
	.full(fullProc33West),
	.dataIn(dataOutProc33West),
	.rd(rdProc32East),
	.empty(emptyProc32East),
	.dataOut(dataInProc32East));
	
	//FIFO 32 TO 33
fifo fifo_proc32_to_proc33(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc32East),
	.full(fullProc32East),
	.dataIn(dataOutProc32East),
	.rd(rdProc33West),
	.empty(emptyProc33West),
	.dataOut(dataInProc33West));
	
	//FIFO 33 TO 20 
fifo fifo_proc33_to_proc20(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc33North),
	.full(fullProc33North),
	.dataIn(dataOutProc33North),
	.rd(rdProc20South),
	.empty(emptyProc20South),
	.dataOut(dataInProc20South));
	
	//FIFO 20 TO 33
fifo fifo_proc20_to_proc33(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc20South),
	.full(fullProc20South),
	.dataIn(dataOutProc20South),
	.rd(rdProc33North),
	.empty(emptyProc33North),
	.dataOut(dataInProc33North));

	//FIFO 34 TO 33 
fifo fifo_proc34_to_proc33(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc34West),
	.full(fullProc34West),
	.dataIn(dataOutProc34West),
	.rd(rdProc33East),
	.empty(emptyProc33East),
	.dataOut(dataInProc33East));
	
	//FIFO 33 TO 34
fifo fifo_proc33_to_proc34(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc33East),
	.full(fullProc33East),
	.dataIn(dataOutProc33East),
	.rd(rdProc34West),
	.empty(emptyProc34West),
	.dataOut(dataInProc34West));
	
	//FIFO 34 TO 21 
fifo fifo_proc34_to_proc21(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc34North),
	.full(fullProc34North),
	.dataIn(dataOutProc34North),
	.rd(rdProc21South),
	.empty(emptyProc21South),
	.dataOut(dataInProc21South));
	
	//FIFO 21 TO 34
fifo fifo_proc21_to_proc34(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc21South),
	.full(fullProc21South),
	.dataIn(dataOutProc21South),
	.rd(rdProc34North),
	.empty(emptyProc34North),
	.dataOut(dataInProc34North));

	//FIFO 35 TO 34 
fifo fifo_proc35_to_proc34(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc35West),
	.full(fullProc35West),
	.dataIn(dataOutProc35West),
	.rd(rdProc34East),
	.empty(emptyProc34East),
	.dataOut(dataInProc34East));
	
	//FIFO 34 TO 35
fifo fifo_proc34_to_proc35(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc34East),
	.full(fullProc34East),
	.dataIn(dataOutProc34East),
	.rd(rdProc35West),
	.empty(emptyProc35West),
	.dataOut(dataInProc35West));
	
	//FIFO 35 TO 22 
fifo fifo_proc35_to_proc22(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc35North),
	.full(fullProc35North),
	.dataIn(dataOutProc35North),
	.rd(rdProc22South),
	.empty(emptyProc22South),
	.dataOut(dataInProc22South));
	
	//FIFO 22 TO 35
fifo fifo_proc22_to_proc35(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc22South),
	.full(fullProc22South),
	.dataIn(dataOutProc22South),
	.rd(rdProc35North),
	.empty(emptyProc35North),
	.dataOut(dataInProc35North));

	//FIFO 36 TO 35 
fifo fifo_proc36_to_proc35(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc36West),
	.full(fullProc36West),
	.dataIn(dataOutProc36West),
	.rd(rdProc35East),
	.empty(emptyProc35East),
	.dataOut(dataInProc35East));
	
	//FIFO 35 TO 36
fifo fifo_proc35_to_proc36(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc35East),
	.full(fullProc35East),
	.dataIn(dataOutProc35East),
	.rd(rdProc36West),
	.empty(emptyProc36West),
	.dataOut(dataInProc36West));
	
	//FIFO 36 TO 23 
fifo fifo_proc36_to_proc23(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc36North),
	.full(fullProc36North),
	.dataIn(dataOutProc36North),
	.rd(rdProc23South),
	.empty(emptyProc23South),
	.dataOut(dataInProc23South));
	
	//FIFO 23 TO 36
fifo fifo_proc23_to_proc36(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc23South),
	.full(fullProc23South),
	.dataIn(dataOutProc23South),
	.rd(rdProc36North),
	.empty(emptyProc36North),
	.dataOut(dataInProc36North));

	//FIFO 37 TO 36 
fifo fifo_proc37_to_proc36(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc37West),
	.full(fullProc37West),
	.dataIn(dataOutProc37West),
	.rd(rdProc36East),
	.empty(emptyProc36East),
	.dataOut(dataInProc36East));
	
	//FIFO 36 TO 37
fifo fifo_proc36_to_proc37(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc36East),
	.full(fullProc36East),
	.dataIn(dataOutProc36East),
	.rd(rdProc37West),
	.empty(emptyProc37West),
	.dataOut(dataInProc37West));
	
	//FIFO 37 TO 24 
fifo fifo_proc37_to_proc24(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc37North),
	.full(fullProc37North),
	.dataIn(dataOutProc37North),
	.rd(rdProc24South),
	.empty(emptyProc24South),
	.dataOut(dataInProc24South));
	
	//FIFO 24 TO 37
fifo fifo_proc24_to_proc37(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc24South),
	.full(fullProc24South),
	.dataIn(dataOutProc24South),
	.rd(rdProc37North),
	.empty(emptyProc37North),
	.dataOut(dataInProc37North));

	//FIFO 38 TO 37 
fifo fifo_proc38_to_proc37(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc38West),
	.full(fullProc38West),
	.dataIn(dataOutProc38West),
	.rd(rdProc37East),
	.empty(emptyProc37East),
	.dataOut(dataInProc37East));
	
	//FIFO 37 TO 38
fifo fifo_proc37_to_proc38(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc37East),
	.full(fullProc37East),
	.dataIn(dataOutProc37East),
	.rd(rdProc38West),
	.empty(emptyProc38West),
	.dataOut(dataInProc38West));
	
	//FIFO 38 TO 25 
fifo fifo_proc38_to_proc25(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc38North),
	.full(fullProc38North),
	.dataIn(dataOutProc38North),
	.rd(rdProc25South),
	.empty(emptyProc25South),
	.dataOut(dataInProc25South));
	
	//FIFO 25 TO 38
fifo fifo_proc25_to_proc38(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc25South),
	.full(fullProc25South),
	.dataIn(dataOutProc25South),
	.rd(rdProc38North),
	.empty(emptyProc38North),
	.dataOut(dataInProc38North));

	//FIFO 39 TO 26 
fifo fifo_proc39_to_proc26(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc39North),
	.full(fullProc39North),
	.dataIn(dataOutProc39North),
	.rd(rdProc26South),
	.empty(emptyProc26South),
	.dataOut(dataInProc26South));
	
	//FIFO 26 TO 39
fifo fifo_proc26_to_proc39(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc26South),
	.full(fullProc26South),
	.dataIn(dataOutProc26South),
	.rd(rdProc39North),
	.empty(emptyProc39North),
	.dataOut(dataInProc39North));

	//FIFO 40 TO 39 
fifo fifo_proc40_to_proc39(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc40West),
	.full(fullProc40West),
	.dataIn(dataOutProc40West),
	.rd(rdProc39East),
	.empty(emptyProc39East),
	.dataOut(dataInProc39East));
	
	//FIFO 39 TO 40
fifo fifo_proc39_to_proc40(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc39East),
	.full(fullProc39East),
	.dataIn(dataOutProc39East),
	.rd(rdProc40West),
	.empty(emptyProc40West),
	.dataOut(dataInProc40West));
	
	//FIFO 40 TO 27 
fifo fifo_proc40_to_proc27(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc40North),
	.full(fullProc40North),
	.dataIn(dataOutProc40North),
	.rd(rdProc27South),
	.empty(emptyProc27South),
	.dataOut(dataInProc27South));
	
	//FIFO 27 TO 40
fifo fifo_proc27_to_proc40(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc27South),
	.full(fullProc27South),
	.dataIn(dataOutProc27South),
	.rd(rdProc40North),
	.empty(emptyProc40North),
	.dataOut(dataInProc40North));

	//FIFO 41 TO 40 
fifo fifo_proc41_to_proc40(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc41West),
	.full(fullProc41West),
	.dataIn(dataOutProc41West),
	.rd(rdProc40East),
	.empty(emptyProc40East),
	.dataOut(dataInProc40East));
	
	//FIFO 40 TO 41
fifo fifo_proc40_to_proc41(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc40East),
	.full(fullProc40East),
	.dataIn(dataOutProc40East),
	.rd(rdProc41West),
	.empty(emptyProc41West),
	.dataOut(dataInProc41West));
	
	//FIFO 41 TO 28 
fifo fifo_proc41_to_proc28(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc41North),
	.full(fullProc41North),
	.dataIn(dataOutProc41North),
	.rd(rdProc28South),
	.empty(emptyProc28South),
	.dataOut(dataInProc28South));
	
	//FIFO 28 TO 41
fifo fifo_proc28_to_proc41(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc28South),
	.full(fullProc28South),
	.dataIn(dataOutProc28South),
	.rd(rdProc41North),
	.empty(emptyProc41North),
	.dataOut(dataInProc41North));

	//FIFO 42 TO 41 
fifo fifo_proc42_to_proc41(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc42West),
	.full(fullProc42West),
	.dataIn(dataOutProc42West),
	.rd(rdProc41East),
	.empty(emptyProc41East),
	.dataOut(dataInProc41East));
	
	//FIFO 41 TO 42
fifo fifo_proc41_to_proc42(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc41East),
	.full(fullProc41East),
	.dataIn(dataOutProc41East),
	.rd(rdProc42West),
	.empty(emptyProc42West),
	.dataOut(dataInProc42West));
	
	//FIFO 42 TO 29 
fifo fifo_proc42_to_proc29(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc42North),
	.full(fullProc42North),
	.dataIn(dataOutProc42North),
	.rd(rdProc29South),
	.empty(emptyProc29South),
	.dataOut(dataInProc29South));
	
	//FIFO 29 TO 42
fifo fifo_proc29_to_proc42(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc29South),
	.full(fullProc29South),
	.dataIn(dataOutProc29South),
	.rd(rdProc42North),
	.empty(emptyProc42North),
	.dataOut(dataInProc42North));

	//FIFO 43 TO 42 
fifo fifo_proc43_to_proc42(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc43West),
	.full(fullProc43West),
	.dataIn(dataOutProc43West),
	.rd(rdProc42East),
	.empty(emptyProc42East),
	.dataOut(dataInProc42East));
	
	//FIFO 42 TO 43
fifo fifo_proc42_to_proc43(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc42East),
	.full(fullProc42East),
	.dataIn(dataOutProc42East),
	.rd(rdProc43West),
	.empty(emptyProc43West),
	.dataOut(dataInProc43West));
	
	//FIFO 43 TO 30 
fifo fifo_proc43_to_proc30(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc43North),
	.full(fullProc43North),
	.dataIn(dataOutProc43North),
	.rd(rdProc30South),
	.empty(emptyProc30South),
	.dataOut(dataInProc30South));
	
	//FIFO 30 TO 43
fifo fifo_proc30_to_proc43(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc30South),
	.full(fullProc30South),
	.dataIn(dataOutProc30South),
	.rd(rdProc43North),
	.empty(emptyProc43North),
	.dataOut(dataInProc43North));

	//FIFO 44 TO 43 
fifo fifo_proc44_to_proc43(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc44West),
	.full(fullProc44West),
	.dataIn(dataOutProc44West),
	.rd(rdProc43East),
	.empty(emptyProc43East),
	.dataOut(dataInProc43East));
	
	//FIFO 43 TO 44
fifo fifo_proc43_to_proc44(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc43East),
	.full(fullProc43East),
	.dataIn(dataOutProc43East),
	.rd(rdProc44West),
	.empty(emptyProc44West),
	.dataOut(dataInProc44West));
	
	//FIFO 44 TO 31 
fifo fifo_proc44_to_proc31(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc44North),
	.full(fullProc44North),
	.dataIn(dataOutProc44North),
	.rd(rdProc31South),
	.empty(emptyProc31South),
	.dataOut(dataInProc31South));
	
	//FIFO 31 TO 44
fifo fifo_proc31_to_proc44(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc31South),
	.full(fullProc31South),
	.dataIn(dataOutProc31South),
	.rd(rdProc44North),
	.empty(emptyProc44North),
	.dataOut(dataInProc44North));

	//FIFO 45 TO 44 
fifo fifo_proc45_to_proc44(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc45West),
	.full(fullProc45West),
	.dataIn(dataOutProc45West),
	.rd(rdProc44East),
	.empty(emptyProc44East),
	.dataOut(dataInProc44East));
	
	//FIFO 44 TO 45
fifo fifo_proc44_to_proc45(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc44East),
	.full(fullProc44East),
	.dataIn(dataOutProc44East),
	.rd(rdProc45West),
	.empty(emptyProc45West),
	.dataOut(dataInProc45West));
	
	//FIFO 45 TO 32 
fifo fifo_proc45_to_proc32(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc45North),
	.full(fullProc45North),
	.dataIn(dataOutProc45North),
	.rd(rdProc32South),
	.empty(emptyProc32South),
	.dataOut(dataInProc32South));
	
	//FIFO 32 TO 45
fifo fifo_proc32_to_proc45(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc32South),
	.full(fullProc32South),
	.dataIn(dataOutProc32South),
	.rd(rdProc45North),
	.empty(emptyProc45North),
	.dataOut(dataInProc45North));

	//FIFO 46 TO 45 
fifo fifo_proc46_to_proc45(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc46West),
	.full(fullProc46West),
	.dataIn(dataOutProc46West),
	.rd(rdProc45East),
	.empty(emptyProc45East),
	.dataOut(dataInProc45East));
	
	//FIFO 45 TO 46
fifo fifo_proc45_to_proc46(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc45East),
	.full(fullProc45East),
	.dataIn(dataOutProc45East),
	.rd(rdProc46West),
	.empty(emptyProc46West),
	.dataOut(dataInProc46West));
	
	//FIFO 46 TO 33 
fifo fifo_proc46_to_proc33(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc46North),
	.full(fullProc46North),
	.dataIn(dataOutProc46North),
	.rd(rdProc33South),
	.empty(emptyProc33South),
	.dataOut(dataInProc33South));
	
	//FIFO 33 TO 46
fifo fifo_proc33_to_proc46(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc33South),
	.full(fullProc33South),
	.dataIn(dataOutProc33South),
	.rd(rdProc46North),
	.empty(emptyProc46North),
	.dataOut(dataInProc46North));

	//FIFO 47 TO 46 
fifo fifo_proc47_to_proc46(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc47West),
	.full(fullProc47West),
	.dataIn(dataOutProc47West),
	.rd(rdProc46East),
	.empty(emptyProc46East),
	.dataOut(dataInProc46East));
	
	//FIFO 46 TO 47
fifo fifo_proc46_to_proc47(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc46East),
	.full(fullProc46East),
	.dataIn(dataOutProc46East),
	.rd(rdProc47West),
	.empty(emptyProc47West),
	.dataOut(dataInProc47West));
	
	//FIFO 47 TO 34 
fifo fifo_proc47_to_proc34(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc47North),
	.full(fullProc47North),
	.dataIn(dataOutProc47North),
	.rd(rdProc34South),
	.empty(emptyProc34South),
	.dataOut(dataInProc34South));
	
	//FIFO 34 TO 47
fifo fifo_proc34_to_proc47(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc34South),
	.full(fullProc34South),
	.dataIn(dataOutProc34South),
	.rd(rdProc47North),
	.empty(emptyProc47North),
	.dataOut(dataInProc47North));

	//FIFO 48 TO 47 
fifo fifo_proc48_to_proc47(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc48West),
	.full(fullProc48West),
	.dataIn(dataOutProc48West),
	.rd(rdProc47East),
	.empty(emptyProc47East),
	.dataOut(dataInProc47East));
	
	//FIFO 47 TO 48
fifo fifo_proc47_to_proc48(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc47East),
	.full(fullProc47East),
	.dataIn(dataOutProc47East),
	.rd(rdProc48West),
	.empty(emptyProc48West),
	.dataOut(dataInProc48West));
	
	//FIFO 48 TO 35 
fifo fifo_proc48_to_proc35(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc48North),
	.full(fullProc48North),
	.dataIn(dataOutProc48North),
	.rd(rdProc35South),
	.empty(emptyProc35South),
	.dataOut(dataInProc35South));
	
	//FIFO 35 TO 48
fifo fifo_proc35_to_proc48(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc35South),
	.full(fullProc35South),
	.dataIn(dataOutProc35South),
	.rd(rdProc48North),
	.empty(emptyProc48North),
	.dataOut(dataInProc48North));

	//FIFO 49 TO 48 
fifo fifo_proc49_to_proc48(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc49West),
	.full(fullProc49West),
	.dataIn(dataOutProc49West),
	.rd(rdProc48East),
	.empty(emptyProc48East),
	.dataOut(dataInProc48East));
	
	//FIFO 48 TO 49
fifo fifo_proc48_to_proc49(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc48East),
	.full(fullProc48East),
	.dataIn(dataOutProc48East),
	.rd(rdProc49West),
	.empty(emptyProc49West),
	.dataOut(dataInProc49West));
	
	//FIFO 49 TO 36 
fifo fifo_proc49_to_proc36(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc49North),
	.full(fullProc49North),
	.dataIn(dataOutProc49North),
	.rd(rdProc36South),
	.empty(emptyProc36South),
	.dataOut(dataInProc36South));
	
	//FIFO 36 TO 49
fifo fifo_proc36_to_proc49(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc36South),
	.full(fullProc36South),
	.dataIn(dataOutProc36South),
	.rd(rdProc49North),
	.empty(emptyProc49North),
	.dataOut(dataInProc49North));

	//FIFO 50 TO 49 
fifo fifo_proc50_to_proc49(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc50West),
	.full(fullProc50West),
	.dataIn(dataOutProc50West),
	.rd(rdProc49East),
	.empty(emptyProc49East),
	.dataOut(dataInProc49East));
	
	//FIFO 49 TO 50
fifo fifo_proc49_to_proc50(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc49East),
	.full(fullProc49East),
	.dataIn(dataOutProc49East),
	.rd(rdProc50West),
	.empty(emptyProc50West),
	.dataOut(dataInProc50West));
	
	//FIFO 50 TO 37 
fifo fifo_proc50_to_proc37(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc50North),
	.full(fullProc50North),
	.dataIn(dataOutProc50North),
	.rd(rdProc37South),
	.empty(emptyProc37South),
	.dataOut(dataInProc37South));
	
	//FIFO 37 TO 50
fifo fifo_proc37_to_proc50(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc37South),
	.full(fullProc37South),
	.dataIn(dataOutProc37South),
	.rd(rdProc50North),
	.empty(emptyProc50North),
	.dataOut(dataInProc50North));

	//FIFO 51 TO 50 
fifo fifo_proc51_to_proc50(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc51West),
	.full(fullProc51West),
	.dataIn(dataOutProc51West),
	.rd(rdProc50East),
	.empty(emptyProc50East),
	.dataOut(dataInProc50East));
	
	//FIFO 50 TO 51
fifo fifo_proc50_to_proc51(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc50East),
	.full(fullProc50East),
	.dataIn(dataOutProc50East),
	.rd(rdProc51West),
	.empty(emptyProc51West),
	.dataOut(dataInProc51West));
	
	//FIFO 51 TO 38 
fifo fifo_proc51_to_proc38(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc51North),
	.full(fullProc51North),
	.dataIn(dataOutProc51North),
	.rd(rdProc38South),
	.empty(emptyProc38South),
	.dataOut(dataInProc38South));
	
	//FIFO 38 TO 51
fifo fifo_proc38_to_proc51(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc38South),
	.full(fullProc38South),
	.dataIn(dataOutProc38South),
	.rd(rdProc51North),
	.empty(emptyProc51North),
	.dataOut(dataInProc51North));

	//FIFO 52 TO 39 
fifo fifo_proc52_to_proc39(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc52North),
	.full(fullProc52North),
	.dataIn(dataOutProc52North),
	.rd(rdProc39South),
	.empty(emptyProc39South),
	.dataOut(dataInProc39South));
	
	//FIFO 39 TO 52
fifo fifo_proc39_to_proc52(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc39South),
	.full(fullProc39South),
	.dataIn(dataOutProc39South),
	.rd(rdProc52North),
	.empty(emptyProc52North),
	.dataOut(dataInProc52North));

	//FIFO 53 TO 52 
fifo fifo_proc53_to_proc52(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc53West),
	.full(fullProc53West),
	.dataIn(dataOutProc53West),
	.rd(rdProc52East),
	.empty(emptyProc52East),
	.dataOut(dataInProc52East));
	
	//FIFO 52 TO 53
fifo fifo_proc52_to_proc53(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc52East),
	.full(fullProc52East),
	.dataIn(dataOutProc52East),
	.rd(rdProc53West),
	.empty(emptyProc53West),
	.dataOut(dataInProc53West));
	
	//FIFO 53 TO 40 
fifo fifo_proc53_to_proc40(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc53North),
	.full(fullProc53North),
	.dataIn(dataOutProc53North),
	.rd(rdProc40South),
	.empty(emptyProc40South),
	.dataOut(dataInProc40South));
	
	//FIFO 40 TO 53
fifo fifo_proc40_to_proc53(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc40South),
	.full(fullProc40South),
	.dataIn(dataOutProc40South),
	.rd(rdProc53North),
	.empty(emptyProc53North),
	.dataOut(dataInProc53North));

	//FIFO 54 TO 53 
fifo fifo_proc54_to_proc53(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc54West),
	.full(fullProc54West),
	.dataIn(dataOutProc54West),
	.rd(rdProc53East),
	.empty(emptyProc53East),
	.dataOut(dataInProc53East));
	
	//FIFO 53 TO 54
fifo fifo_proc53_to_proc54(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc53East),
	.full(fullProc53East),
	.dataIn(dataOutProc53East),
	.rd(rdProc54West),
	.empty(emptyProc54West),
	.dataOut(dataInProc54West));
	
	//FIFO 54 TO 41 
fifo fifo_proc54_to_proc41(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc54North),
	.full(fullProc54North),
	.dataIn(dataOutProc54North),
	.rd(rdProc41South),
	.empty(emptyProc41South),
	.dataOut(dataInProc41South));
	
	//FIFO 41 TO 54
fifo fifo_proc41_to_proc54(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc41South),
	.full(fullProc41South),
	.dataIn(dataOutProc41South),
	.rd(rdProc54North),
	.empty(emptyProc54North),
	.dataOut(dataInProc54North));

	//FIFO 55 TO 54 
fifo fifo_proc55_to_proc54(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc55West),
	.full(fullProc55West),
	.dataIn(dataOutProc55West),
	.rd(rdProc54East),
	.empty(emptyProc54East),
	.dataOut(dataInProc54East));
	
	//FIFO 54 TO 55
fifo fifo_proc54_to_proc55(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc54East),
	.full(fullProc54East),
	.dataIn(dataOutProc54East),
	.rd(rdProc55West),
	.empty(emptyProc55West),
	.dataOut(dataInProc55West));
	
	//FIFO 55 TO 42 
fifo fifo_proc55_to_proc42(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc55North),
	.full(fullProc55North),
	.dataIn(dataOutProc55North),
	.rd(rdProc42South),
	.empty(emptyProc42South),
	.dataOut(dataInProc42South));
	
	//FIFO 42 TO 55
fifo fifo_proc42_to_proc55(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc42South),
	.full(fullProc42South),
	.dataIn(dataOutProc42South),
	.rd(rdProc55North),
	.empty(emptyProc55North),
	.dataOut(dataInProc55North));

	//FIFO 56 TO 55 
fifo fifo_proc56_to_proc55(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc56West),
	.full(fullProc56West),
	.dataIn(dataOutProc56West),
	.rd(rdProc55East),
	.empty(emptyProc55East),
	.dataOut(dataInProc55East));
	
	//FIFO 55 TO 56
fifo fifo_proc55_to_proc56(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc55East),
	.full(fullProc55East),
	.dataIn(dataOutProc55East),
	.rd(rdProc56West),
	.empty(emptyProc56West),
	.dataOut(dataInProc56West));
	
	//FIFO 56 TO 43 
fifo fifo_proc56_to_proc43(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc56North),
	.full(fullProc56North),
	.dataIn(dataOutProc56North),
	.rd(rdProc43South),
	.empty(emptyProc43South),
	.dataOut(dataInProc43South));
	
	//FIFO 43 TO 56
fifo fifo_proc43_to_proc56(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc43South),
	.full(fullProc43South),
	.dataIn(dataOutProc43South),
	.rd(rdProc56North),
	.empty(emptyProc56North),
	.dataOut(dataInProc56North));

	//FIFO 57 TO 56 
fifo fifo_proc57_to_proc56(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc57West),
	.full(fullProc57West),
	.dataIn(dataOutProc57West),
	.rd(rdProc56East),
	.empty(emptyProc56East),
	.dataOut(dataInProc56East));
	
	//FIFO 56 TO 57
fifo fifo_proc56_to_proc57(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc56East),
	.full(fullProc56East),
	.dataIn(dataOutProc56East),
	.rd(rdProc57West),
	.empty(emptyProc57West),
	.dataOut(dataInProc57West));
	
	//FIFO 57 TO 44 
fifo fifo_proc57_to_proc44(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc57North),
	.full(fullProc57North),
	.dataIn(dataOutProc57North),
	.rd(rdProc44South),
	.empty(emptyProc44South),
	.dataOut(dataInProc44South));
	
	//FIFO 44 TO 57
fifo fifo_proc44_to_proc57(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc44South),
	.full(fullProc44South),
	.dataIn(dataOutProc44South),
	.rd(rdProc57North),
	.empty(emptyProc57North),
	.dataOut(dataInProc57North));

	//FIFO 58 TO 57 
fifo fifo_proc58_to_proc57(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc58West),
	.full(fullProc58West),
	.dataIn(dataOutProc58West),
	.rd(rdProc57East),
	.empty(emptyProc57East),
	.dataOut(dataInProc57East));
	
	//FIFO 57 TO 58
fifo fifo_proc57_to_proc58(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc57East),
	.full(fullProc57East),
	.dataIn(dataOutProc57East),
	.rd(rdProc58West),
	.empty(emptyProc58West),
	.dataOut(dataInProc58West));
	
	//FIFO 58 TO 45 
fifo fifo_proc58_to_proc45(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc58North),
	.full(fullProc58North),
	.dataIn(dataOutProc58North),
	.rd(rdProc45South),
	.empty(emptyProc45South),
	.dataOut(dataInProc45South));
	
	//FIFO 45 TO 58
fifo fifo_proc45_to_proc58(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc45South),
	.full(fullProc45South),
	.dataIn(dataOutProc45South),
	.rd(rdProc58North),
	.empty(emptyProc58North),
	.dataOut(dataInProc58North));

	//FIFO 59 TO 58 
fifo fifo_proc59_to_proc58(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc59West),
	.full(fullProc59West),
	.dataIn(dataOutProc59West),
	.rd(rdProc58East),
	.empty(emptyProc58East),
	.dataOut(dataInProc58East));
	
	//FIFO 58 TO 59
fifo fifo_proc58_to_proc59(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc58East),
	.full(fullProc58East),
	.dataIn(dataOutProc58East),
	.rd(rdProc59West),
	.empty(emptyProc59West),
	.dataOut(dataInProc59West));
	
	//FIFO 59 TO 46 
fifo fifo_proc59_to_proc46(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc59North),
	.full(fullProc59North),
	.dataIn(dataOutProc59North),
	.rd(rdProc46South),
	.empty(emptyProc46South),
	.dataOut(dataInProc46South));
	
	//FIFO 46 TO 59
fifo fifo_proc46_to_proc59(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc46South),
	.full(fullProc46South),
	.dataIn(dataOutProc46South),
	.rd(rdProc59North),
	.empty(emptyProc59North),
	.dataOut(dataInProc59North));

	//FIFO 60 TO 59 
fifo fifo_proc60_to_proc59(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc60West),
	.full(fullProc60West),
	.dataIn(dataOutProc60West),
	.rd(rdProc59East),
	.empty(emptyProc59East),
	.dataOut(dataInProc59East));
	
	//FIFO 59 TO 60
fifo fifo_proc59_to_proc60(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc59East),
	.full(fullProc59East),
	.dataIn(dataOutProc59East),
	.rd(rdProc60West),
	.empty(emptyProc60West),
	.dataOut(dataInProc60West));
	
	//FIFO 60 TO 47 
fifo fifo_proc60_to_proc47(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc60North),
	.full(fullProc60North),
	.dataIn(dataOutProc60North),
	.rd(rdProc47South),
	.empty(emptyProc47South),
	.dataOut(dataInProc47South));
	
	//FIFO 47 TO 60
fifo fifo_proc47_to_proc60(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc47South),
	.full(fullProc47South),
	.dataIn(dataOutProc47South),
	.rd(rdProc60North),
	.empty(emptyProc60North),
	.dataOut(dataInProc60North));

	//FIFO 61 TO 60 
fifo fifo_proc61_to_proc60(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc61West),
	.full(fullProc61West),
	.dataIn(dataOutProc61West),
	.rd(rdProc60East),
	.empty(emptyProc60East),
	.dataOut(dataInProc60East));
	
	//FIFO 60 TO 61
fifo fifo_proc60_to_proc61(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc60East),
	.full(fullProc60East),
	.dataIn(dataOutProc60East),
	.rd(rdProc61West),
	.empty(emptyProc61West),
	.dataOut(dataInProc61West));
	
	//FIFO 61 TO 48 
fifo fifo_proc61_to_proc48(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc61North),
	.full(fullProc61North),
	.dataIn(dataOutProc61North),
	.rd(rdProc48South),
	.empty(emptyProc48South),
	.dataOut(dataInProc48South));
	
	//FIFO 48 TO 61
fifo fifo_proc48_to_proc61(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc48South),
	.full(fullProc48South),
	.dataIn(dataOutProc48South),
	.rd(rdProc61North),
	.empty(emptyProc61North),
	.dataOut(dataInProc61North));

	//FIFO 62 TO 61 
fifo fifo_proc62_to_proc61(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc62West),
	.full(fullProc62West),
	.dataIn(dataOutProc62West),
	.rd(rdProc61East),
	.empty(emptyProc61East),
	.dataOut(dataInProc61East));
	
	//FIFO 61 TO 62
fifo fifo_proc61_to_proc62(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc61East),
	.full(fullProc61East),
	.dataIn(dataOutProc61East),
	.rd(rdProc62West),
	.empty(emptyProc62West),
	.dataOut(dataInProc62West));
	
	//FIFO 62 TO 49 
fifo fifo_proc62_to_proc49(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc62North),
	.full(fullProc62North),
	.dataIn(dataOutProc62North),
	.rd(rdProc49South),
	.empty(emptyProc49South),
	.dataOut(dataInProc49South));
	
	//FIFO 49 TO 62
fifo fifo_proc49_to_proc62(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc49South),
	.full(fullProc49South),
	.dataIn(dataOutProc49South),
	.rd(rdProc62North),
	.empty(emptyProc62North),
	.dataOut(dataInProc62North));

	//FIFO 63 TO 62 
fifo fifo_proc63_to_proc62(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc63West),
	.full(fullProc63West),
	.dataIn(dataOutProc63West),
	.rd(rdProc62East),
	.empty(emptyProc62East),
	.dataOut(dataInProc62East));
	
	//FIFO 62 TO 63
fifo fifo_proc62_to_proc63(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc62East),
	.full(fullProc62East),
	.dataIn(dataOutProc62East),
	.rd(rdProc63West),
	.empty(emptyProc63West),
	.dataOut(dataInProc63West));
	
	//FIFO 63 TO 50 
fifo fifo_proc63_to_proc50(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc63North),
	.full(fullProc63North),
	.dataIn(dataOutProc63North),
	.rd(rdProc50South),
	.empty(emptyProc50South),
	.dataOut(dataInProc50South));
	
	//FIFO 50 TO 63
fifo fifo_proc50_to_proc63(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc50South),
	.full(fullProc50South),
	.dataIn(dataOutProc50South),
	.rd(rdProc63North),
	.empty(emptyProc63North),
	.dataOut(dataInProc63North));

	//FIFO 64 TO 63 
fifo fifo_proc64_to_proc63(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc64West),
	.full(fullProc64West),
	.dataIn(dataOutProc64West),
	.rd(rdProc63East),
	.empty(emptyProc63East),
	.dataOut(dataInProc63East));
	
	//FIFO 63 TO 64
fifo fifo_proc63_to_proc64(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc63East),
	.full(fullProc63East),
	.dataIn(dataOutProc63East),
	.rd(rdProc64West),
	.empty(emptyProc64West),
	.dataOut(dataInProc64West));
	
	//FIFO 64 TO 51 
fifo fifo_proc64_to_proc51(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc64North),
	.full(fullProc64North),
	.dataIn(dataOutProc64North),
	.rd(rdProc51South),
	.empty(emptyProc51South),
	.dataOut(dataInProc51South));
	
	//FIFO 51 TO 64
fifo fifo_proc51_to_proc64(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc51South),
	.full(fullProc51South),
	.dataIn(dataOutProc51South),
	.rd(rdProc64North),
	.empty(emptyProc64North),
	.dataOut(dataInProc64North));

	//FIFO 65 TO 52 
fifo fifo_proc65_to_proc52(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc65North),
	.full(fullProc65North),
	.dataIn(dataOutProc65North),
	.rd(rdProc52South),
	.empty(emptyProc52South),
	.dataOut(dataInProc52South));
	
	//FIFO 52 TO 65
fifo fifo_proc52_to_proc65(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc52South),
	.full(fullProc52South),
	.dataIn(dataOutProc52South),
	.rd(rdProc65North),
	.empty(emptyProc65North),
	.dataOut(dataInProc65North));

	//FIFO 66 TO 65 
fifo fifo_proc66_to_proc65(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc66West),
	.full(fullProc66West),
	.dataIn(dataOutProc66West),
	.rd(rdProc65East),
	.empty(emptyProc65East),
	.dataOut(dataInProc65East));
	
	//FIFO 65 TO 66
fifo fifo_proc65_to_proc66(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc65East),
	.full(fullProc65East),
	.dataIn(dataOutProc65East),
	.rd(rdProc66West),
	.empty(emptyProc66West),
	.dataOut(dataInProc66West));
	
	//FIFO 66 TO 53 
fifo fifo_proc66_to_proc53(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc66North),
	.full(fullProc66North),
	.dataIn(dataOutProc66North),
	.rd(rdProc53South),
	.empty(emptyProc53South),
	.dataOut(dataInProc53South));
	
	//FIFO 53 TO 66
fifo fifo_proc53_to_proc66(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc53South),
	.full(fullProc53South),
	.dataIn(dataOutProc53South),
	.rd(rdProc66North),
	.empty(emptyProc66North),
	.dataOut(dataInProc66North));

	//FIFO 67 TO 66 
fifo fifo_proc67_to_proc66(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc67West),
	.full(fullProc67West),
	.dataIn(dataOutProc67West),
	.rd(rdProc66East),
	.empty(emptyProc66East),
	.dataOut(dataInProc66East));
	
	//FIFO 66 TO 67
fifo fifo_proc66_to_proc67(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc66East),
	.full(fullProc66East),
	.dataIn(dataOutProc66East),
	.rd(rdProc67West),
	.empty(emptyProc67West),
	.dataOut(dataInProc67West));
	
	//FIFO 67 TO 54 
fifo fifo_proc67_to_proc54(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc67North),
	.full(fullProc67North),
	.dataIn(dataOutProc67North),
	.rd(rdProc54South),
	.empty(emptyProc54South),
	.dataOut(dataInProc54South));
	
	//FIFO 54 TO 67
fifo fifo_proc54_to_proc67(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc54South),
	.full(fullProc54South),
	.dataIn(dataOutProc54South),
	.rd(rdProc67North),
	.empty(emptyProc67North),
	.dataOut(dataInProc67North));

	//FIFO 68 TO 67 
fifo fifo_proc68_to_proc67(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc68West),
	.full(fullProc68West),
	.dataIn(dataOutProc68West),
	.rd(rdProc67East),
	.empty(emptyProc67East),
	.dataOut(dataInProc67East));
	
	//FIFO 67 TO 68
fifo fifo_proc67_to_proc68(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc67East),
	.full(fullProc67East),
	.dataIn(dataOutProc67East),
	.rd(rdProc68West),
	.empty(emptyProc68West),
	.dataOut(dataInProc68West));
	
	//FIFO 68 TO 55 
fifo fifo_proc68_to_proc55(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc68North),
	.full(fullProc68North),
	.dataIn(dataOutProc68North),
	.rd(rdProc55South),
	.empty(emptyProc55South),
	.dataOut(dataInProc55South));
	
	//FIFO 55 TO 68
fifo fifo_proc55_to_proc68(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc55South),
	.full(fullProc55South),
	.dataIn(dataOutProc55South),
	.rd(rdProc68North),
	.empty(emptyProc68North),
	.dataOut(dataInProc68North));

	//FIFO 69 TO 68 
fifo fifo_proc69_to_proc68(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc69West),
	.full(fullProc69West),
	.dataIn(dataOutProc69West),
	.rd(rdProc68East),
	.empty(emptyProc68East),
	.dataOut(dataInProc68East));
	
	//FIFO 68 TO 69
fifo fifo_proc68_to_proc69(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc68East),
	.full(fullProc68East),
	.dataIn(dataOutProc68East),
	.rd(rdProc69West),
	.empty(emptyProc69West),
	.dataOut(dataInProc69West));
	
	//FIFO 69 TO 56 
fifo fifo_proc69_to_proc56(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc69North),
	.full(fullProc69North),
	.dataIn(dataOutProc69North),
	.rd(rdProc56South),
	.empty(emptyProc56South),
	.dataOut(dataInProc56South));
	
	//FIFO 56 TO 69
fifo fifo_proc56_to_proc69(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc56South),
	.full(fullProc56South),
	.dataIn(dataOutProc56South),
	.rd(rdProc69North),
	.empty(emptyProc69North),
	.dataOut(dataInProc69North));

	//FIFO 70 TO 69 
fifo fifo_proc70_to_proc69(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc70West),
	.full(fullProc70West),
	.dataIn(dataOutProc70West),
	.rd(rdProc69East),
	.empty(emptyProc69East),
	.dataOut(dataInProc69East));
	
	//FIFO 69 TO 70
fifo fifo_proc69_to_proc70(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc69East),
	.full(fullProc69East),
	.dataIn(dataOutProc69East),
	.rd(rdProc70West),
	.empty(emptyProc70West),
	.dataOut(dataInProc70West));
	
	//FIFO 70 TO 57 
fifo fifo_proc70_to_proc57(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc70North),
	.full(fullProc70North),
	.dataIn(dataOutProc70North),
	.rd(rdProc57South),
	.empty(emptyProc57South),
	.dataOut(dataInProc57South));
	
	//FIFO 57 TO 70
fifo fifo_proc57_to_proc70(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc57South),
	.full(fullProc57South),
	.dataIn(dataOutProc57South),
	.rd(rdProc70North),
	.empty(emptyProc70North),
	.dataOut(dataInProc70North));

	//FIFO 71 TO 70 
fifo fifo_proc71_to_proc70(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc71West),
	.full(fullProc71West),
	.dataIn(dataOutProc71West),
	.rd(rdProc70East),
	.empty(emptyProc70East),
	.dataOut(dataInProc70East));
	
	//FIFO 70 TO 71
fifo fifo_proc70_to_proc71(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc70East),
	.full(fullProc70East),
	.dataIn(dataOutProc70East),
	.rd(rdProc71West),
	.empty(emptyProc71West),
	.dataOut(dataInProc71West));
	
	//FIFO 71 TO 58 
fifo fifo_proc71_to_proc58(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc71North),
	.full(fullProc71North),
	.dataIn(dataOutProc71North),
	.rd(rdProc58South),
	.empty(emptyProc58South),
	.dataOut(dataInProc58South));
	
	//FIFO 58 TO 71
fifo fifo_proc58_to_proc71(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc58South),
	.full(fullProc58South),
	.dataIn(dataOutProc58South),
	.rd(rdProc71North),
	.empty(emptyProc71North),
	.dataOut(dataInProc71North));

	//FIFO 72 TO 71 
fifo fifo_proc72_to_proc71(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc72West),
	.full(fullProc72West),
	.dataIn(dataOutProc72West),
	.rd(rdProc71East),
	.empty(emptyProc71East),
	.dataOut(dataInProc71East));
	
	//FIFO 71 TO 72
fifo fifo_proc71_to_proc72(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc71East),
	.full(fullProc71East),
	.dataIn(dataOutProc71East),
	.rd(rdProc72West),
	.empty(emptyProc72West),
	.dataOut(dataInProc72West));
	
	//FIFO 72 TO 59 
fifo fifo_proc72_to_proc59(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc72North),
	.full(fullProc72North),
	.dataIn(dataOutProc72North),
	.rd(rdProc59South),
	.empty(emptyProc59South),
	.dataOut(dataInProc59South));
	
	//FIFO 59 TO 72
fifo fifo_proc59_to_proc72(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc59South),
	.full(fullProc59South),
	.dataIn(dataOutProc59South),
	.rd(rdProc72North),
	.empty(emptyProc72North),
	.dataOut(dataInProc72North));

	//FIFO 73 TO 72 
fifo fifo_proc73_to_proc72(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc73West),
	.full(fullProc73West),
	.dataIn(dataOutProc73West),
	.rd(rdProc72East),
	.empty(emptyProc72East),
	.dataOut(dataInProc72East));
	
	//FIFO 72 TO 73
fifo fifo_proc72_to_proc73(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc72East),
	.full(fullProc72East),
	.dataIn(dataOutProc72East),
	.rd(rdProc73West),
	.empty(emptyProc73West),
	.dataOut(dataInProc73West));
	
	//FIFO 73 TO 60 
fifo fifo_proc73_to_proc60(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc73North),
	.full(fullProc73North),
	.dataIn(dataOutProc73North),
	.rd(rdProc60South),
	.empty(emptyProc60South),
	.dataOut(dataInProc60South));
	
	//FIFO 60 TO 73
fifo fifo_proc60_to_proc73(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc60South),
	.full(fullProc60South),
	.dataIn(dataOutProc60South),
	.rd(rdProc73North),
	.empty(emptyProc73North),
	.dataOut(dataInProc73North));

	//FIFO 74 TO 73 
fifo fifo_proc74_to_proc73(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc74West),
	.full(fullProc74West),
	.dataIn(dataOutProc74West),
	.rd(rdProc73East),
	.empty(emptyProc73East),
	.dataOut(dataInProc73East));
	
	//FIFO 73 TO 74
fifo fifo_proc73_to_proc74(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc73East),
	.full(fullProc73East),
	.dataIn(dataOutProc73East),
	.rd(rdProc74West),
	.empty(emptyProc74West),
	.dataOut(dataInProc74West));
	
	//FIFO 74 TO 61 
fifo fifo_proc74_to_proc61(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc74North),
	.full(fullProc74North),
	.dataIn(dataOutProc74North),
	.rd(rdProc61South),
	.empty(emptyProc61South),
	.dataOut(dataInProc61South));
	
	//FIFO 61 TO 74
fifo fifo_proc61_to_proc74(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc61South),
	.full(fullProc61South),
	.dataIn(dataOutProc61South),
	.rd(rdProc74North),
	.empty(emptyProc74North),
	.dataOut(dataInProc74North));

	//FIFO 75 TO 74 
fifo fifo_proc75_to_proc74(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc75West),
	.full(fullProc75West),
	.dataIn(dataOutProc75West),
	.rd(rdProc74East),
	.empty(emptyProc74East),
	.dataOut(dataInProc74East));
	
	//FIFO 74 TO 75
fifo fifo_proc74_to_proc75(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc74East),
	.full(fullProc74East),
	.dataIn(dataOutProc74East),
	.rd(rdProc75West),
	.empty(emptyProc75West),
	.dataOut(dataInProc75West));
	
	//FIFO 75 TO 62 
fifo fifo_proc75_to_proc62(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc75North),
	.full(fullProc75North),
	.dataIn(dataOutProc75North),
	.rd(rdProc62South),
	.empty(emptyProc62South),
	.dataOut(dataInProc62South));
	
	//FIFO 62 TO 75
fifo fifo_proc62_to_proc75(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc62South),
	.full(fullProc62South),
	.dataIn(dataOutProc62South),
	.rd(rdProc75North),
	.empty(emptyProc75North),
	.dataOut(dataInProc75North));

	//FIFO 76 TO 75 
fifo fifo_proc76_to_proc75(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc76West),
	.full(fullProc76West),
	.dataIn(dataOutProc76West),
	.rd(rdProc75East),
	.empty(emptyProc75East),
	.dataOut(dataInProc75East));
	
	//FIFO 75 TO 76
fifo fifo_proc75_to_proc76(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc75East),
	.full(fullProc75East),
	.dataIn(dataOutProc75East),
	.rd(rdProc76West),
	.empty(emptyProc76West),
	.dataOut(dataInProc76West));
	
	//FIFO 76 TO 63 
fifo fifo_proc76_to_proc63(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc76North),
	.full(fullProc76North),
	.dataIn(dataOutProc76North),
	.rd(rdProc63South),
	.empty(emptyProc63South),
	.dataOut(dataInProc63South));
	
	//FIFO 63 TO 76
fifo fifo_proc63_to_proc76(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc63South),
	.full(fullProc63South),
	.dataIn(dataOutProc63South),
	.rd(rdProc76North),
	.empty(emptyProc76North),
	.dataOut(dataInProc76North));

	//FIFO 77 TO 76 
fifo fifo_proc77_to_proc76(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc77West),
	.full(fullProc77West),
	.dataIn(dataOutProc77West),
	.rd(rdProc76East),
	.empty(emptyProc76East),
	.dataOut(dataInProc76East));
	
	//FIFO 76 TO 77
fifo fifo_proc76_to_proc77(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc76East),
	.full(fullProc76East),
	.dataIn(dataOutProc76East),
	.rd(rdProc77West),
	.empty(emptyProc77West),
	.dataOut(dataInProc77West));
	
	//FIFO 77 TO 64 
fifo fifo_proc77_to_proc64(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc77North),
	.full(fullProc77North),
	.dataIn(dataOutProc77North),
	.rd(rdProc64South),
	.empty(emptyProc64South),
	.dataOut(dataInProc64South));
	
	//FIFO 64 TO 77
fifo fifo_proc64_to_proc77(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc64South),
	.full(fullProc64South),
	.dataIn(dataOutProc64South),
	.rd(rdProc77North),
	.empty(emptyProc77North),
	.dataOut(dataInProc77North));

	//FIFO 78 TO 65 
fifo fifo_proc78_to_proc65(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc78North),
	.full(fullProc78North),
	.dataIn(dataOutProc78North),
	.rd(rdProc65South),
	.empty(emptyProc65South),
	.dataOut(dataInProc65South));
	
	//FIFO 65 TO 78
fifo fifo_proc65_to_proc78(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc65South),
	.full(fullProc65South),
	.dataIn(dataOutProc65South),
	.rd(rdProc78North),
	.empty(emptyProc78North),
	.dataOut(dataInProc78North));

	//FIFO 79 TO 78 
fifo fifo_proc79_to_proc78(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc79West),
	.full(fullProc79West),
	.dataIn(dataOutProc79West),
	.rd(rdProc78East),
	.empty(emptyProc78East),
	.dataOut(dataInProc78East));
	
	//FIFO 78 TO 79
fifo fifo_proc78_to_proc79(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc78East),
	.full(fullProc78East),
	.dataIn(dataOutProc78East),
	.rd(rdProc79West),
	.empty(emptyProc79West),
	.dataOut(dataInProc79West));
	
	//FIFO 79 TO 66 
fifo fifo_proc79_to_proc66(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc79North),
	.full(fullProc79North),
	.dataIn(dataOutProc79North),
	.rd(rdProc66South),
	.empty(emptyProc66South),
	.dataOut(dataInProc66South));
	
	//FIFO 66 TO 79
fifo fifo_proc66_to_proc79(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc66South),
	.full(fullProc66South),
	.dataIn(dataOutProc66South),
	.rd(rdProc79North),
	.empty(emptyProc79North),
	.dataOut(dataInProc79North));

	//FIFO 80 TO 79 
fifo fifo_proc80_to_proc79(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc80West),
	.full(fullProc80West),
	.dataIn(dataOutProc80West),
	.rd(rdProc79East),
	.empty(emptyProc79East),
	.dataOut(dataInProc79East));
	
	//FIFO 79 TO 80
fifo fifo_proc79_to_proc80(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc79East),
	.full(fullProc79East),
	.dataIn(dataOutProc79East),
	.rd(rdProc80West),
	.empty(emptyProc80West),
	.dataOut(dataInProc80West));
	
	//FIFO 80 TO 67 
fifo fifo_proc80_to_proc67(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc80North),
	.full(fullProc80North),
	.dataIn(dataOutProc80North),
	.rd(rdProc67South),
	.empty(emptyProc67South),
	.dataOut(dataInProc67South));
	
	//FIFO 67 TO 80
fifo fifo_proc67_to_proc80(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc67South),
	.full(fullProc67South),
	.dataIn(dataOutProc67South),
	.rd(rdProc80North),
	.empty(emptyProc80North),
	.dataOut(dataInProc80North));

	//FIFO 81 TO 80 
fifo fifo_proc81_to_proc80(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc81West),
	.full(fullProc81West),
	.dataIn(dataOutProc81West),
	.rd(rdProc80East),
	.empty(emptyProc80East),
	.dataOut(dataInProc80East));
	
	//FIFO 80 TO 81
fifo fifo_proc80_to_proc81(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc80East),
	.full(fullProc80East),
	.dataIn(dataOutProc80East),
	.rd(rdProc81West),
	.empty(emptyProc81West),
	.dataOut(dataInProc81West));
	
	//FIFO 81 TO 68 
fifo fifo_proc81_to_proc68(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc81North),
	.full(fullProc81North),
	.dataIn(dataOutProc81North),
	.rd(rdProc68South),
	.empty(emptyProc68South),
	.dataOut(dataInProc68South));
	
	//FIFO 68 TO 81
fifo fifo_proc68_to_proc81(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc68South),
	.full(fullProc68South),
	.dataIn(dataOutProc68South),
	.rd(rdProc81North),
	.empty(emptyProc81North),
	.dataOut(dataInProc81North));

	//FIFO 82 TO 81 
fifo fifo_proc82_to_proc81(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc82West),
	.full(fullProc82West),
	.dataIn(dataOutProc82West),
	.rd(rdProc81East),
	.empty(emptyProc81East),
	.dataOut(dataInProc81East));
	
	//FIFO 81 TO 82
fifo fifo_proc81_to_proc82(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc81East),
	.full(fullProc81East),
	.dataIn(dataOutProc81East),
	.rd(rdProc82West),
	.empty(emptyProc82West),
	.dataOut(dataInProc82West));
	
	//FIFO 82 TO 69 
fifo fifo_proc82_to_proc69(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc82North),
	.full(fullProc82North),
	.dataIn(dataOutProc82North),
	.rd(rdProc69South),
	.empty(emptyProc69South),
	.dataOut(dataInProc69South));
	
	//FIFO 69 TO 82
fifo fifo_proc69_to_proc82(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc69South),
	.full(fullProc69South),
	.dataIn(dataOutProc69South),
	.rd(rdProc82North),
	.empty(emptyProc82North),
	.dataOut(dataInProc82North));

	//FIFO 83 TO 82 
fifo fifo_proc83_to_proc82(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc83West),
	.full(fullProc83West),
	.dataIn(dataOutProc83West),
	.rd(rdProc82East),
	.empty(emptyProc82East),
	.dataOut(dataInProc82East));
	
	//FIFO 82 TO 83
fifo fifo_proc82_to_proc83(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc82East),
	.full(fullProc82East),
	.dataIn(dataOutProc82East),
	.rd(rdProc83West),
	.empty(emptyProc83West),
	.dataOut(dataInProc83West));
	
	//FIFO 83 TO 70 
fifo fifo_proc83_to_proc70(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc83North),
	.full(fullProc83North),
	.dataIn(dataOutProc83North),
	.rd(rdProc70South),
	.empty(emptyProc70South),
	.dataOut(dataInProc70South));
	
	//FIFO 70 TO 83
fifo fifo_proc70_to_proc83(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc70South),
	.full(fullProc70South),
	.dataIn(dataOutProc70South),
	.rd(rdProc83North),
	.empty(emptyProc83North),
	.dataOut(dataInProc83North));

	//FIFO 84 TO 83 
fifo fifo_proc84_to_proc83(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc84West),
	.full(fullProc84West),
	.dataIn(dataOutProc84West),
	.rd(rdProc83East),
	.empty(emptyProc83East),
	.dataOut(dataInProc83East));
	
	//FIFO 83 TO 84
fifo fifo_proc83_to_proc84(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc83East),
	.full(fullProc83East),
	.dataIn(dataOutProc83East),
	.rd(rdProc84West),
	.empty(emptyProc84West),
	.dataOut(dataInProc84West));
	
	//FIFO 84 TO 71 
fifo fifo_proc84_to_proc71(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc84North),
	.full(fullProc84North),
	.dataIn(dataOutProc84North),
	.rd(rdProc71South),
	.empty(emptyProc71South),
	.dataOut(dataInProc71South));
	
	//FIFO 71 TO 84
fifo fifo_proc71_to_proc84(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc71South),
	.full(fullProc71South),
	.dataIn(dataOutProc71South),
	.rd(rdProc84North),
	.empty(emptyProc84North),
	.dataOut(dataInProc84North));

	//FIFO 85 TO 84 
fifo fifo_proc85_to_proc84(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc85West),
	.full(fullProc85West),
	.dataIn(dataOutProc85West),
	.rd(rdProc84East),
	.empty(emptyProc84East),
	.dataOut(dataInProc84East));
	
	//FIFO 84 TO 85
fifo fifo_proc84_to_proc85(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc84East),
	.full(fullProc84East),
	.dataIn(dataOutProc84East),
	.rd(rdProc85West),
	.empty(emptyProc85West),
	.dataOut(dataInProc85West));
	
	//FIFO 85 TO 72 
fifo fifo_proc85_to_proc72(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc85North),
	.full(fullProc85North),
	.dataIn(dataOutProc85North),
	.rd(rdProc72South),
	.empty(emptyProc72South),
	.dataOut(dataInProc72South));
	
	//FIFO 72 TO 85
fifo fifo_proc72_to_proc85(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc72South),
	.full(fullProc72South),
	.dataIn(dataOutProc72South),
	.rd(rdProc85North),
	.empty(emptyProc85North),
	.dataOut(dataInProc85North));

	//FIFO 86 TO 85 
fifo fifo_proc86_to_proc85(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc86West),
	.full(fullProc86West),
	.dataIn(dataOutProc86West),
	.rd(rdProc85East),
	.empty(emptyProc85East),
	.dataOut(dataInProc85East));
	
	//FIFO 85 TO 86
fifo fifo_proc85_to_proc86(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc85East),
	.full(fullProc85East),
	.dataIn(dataOutProc85East),
	.rd(rdProc86West),
	.empty(emptyProc86West),
	.dataOut(dataInProc86West));
	
	//FIFO 86 TO 73 
fifo fifo_proc86_to_proc73(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc86North),
	.full(fullProc86North),
	.dataIn(dataOutProc86North),
	.rd(rdProc73South),
	.empty(emptyProc73South),
	.dataOut(dataInProc73South));
	
	//FIFO 73 TO 86
fifo fifo_proc73_to_proc86(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc73South),
	.full(fullProc73South),
	.dataIn(dataOutProc73South),
	.rd(rdProc86North),
	.empty(emptyProc86North),
	.dataOut(dataInProc86North));

	//FIFO 87 TO 86 
fifo fifo_proc87_to_proc86(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc87West),
	.full(fullProc87West),
	.dataIn(dataOutProc87West),
	.rd(rdProc86East),
	.empty(emptyProc86East),
	.dataOut(dataInProc86East));
	
	//FIFO 86 TO 87
fifo fifo_proc86_to_proc87(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc86East),
	.full(fullProc86East),
	.dataIn(dataOutProc86East),
	.rd(rdProc87West),
	.empty(emptyProc87West),
	.dataOut(dataInProc87West));
	
	//FIFO 87 TO 74 
fifo fifo_proc87_to_proc74(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc87North),
	.full(fullProc87North),
	.dataIn(dataOutProc87North),
	.rd(rdProc74South),
	.empty(emptyProc74South),
	.dataOut(dataInProc74South));
	
	//FIFO 74 TO 87
fifo fifo_proc74_to_proc87(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc74South),
	.full(fullProc74South),
	.dataIn(dataOutProc74South),
	.rd(rdProc87North),
	.empty(emptyProc87North),
	.dataOut(dataInProc87North));

	//FIFO 88 TO 87 
fifo fifo_proc88_to_proc87(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc88West),
	.full(fullProc88West),
	.dataIn(dataOutProc88West),
	.rd(rdProc87East),
	.empty(emptyProc87East),
	.dataOut(dataInProc87East));
	
	//FIFO 87 TO 88
fifo fifo_proc87_to_proc88(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc87East),
	.full(fullProc87East),
	.dataIn(dataOutProc87East),
	.rd(rdProc88West),
	.empty(emptyProc88West),
	.dataOut(dataInProc88West));
	
	//FIFO 88 TO 75 
fifo fifo_proc88_to_proc75(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc88North),
	.full(fullProc88North),
	.dataIn(dataOutProc88North),
	.rd(rdProc75South),
	.empty(emptyProc75South),
	.dataOut(dataInProc75South));
	
	//FIFO 75 TO 88
fifo fifo_proc75_to_proc88(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc75South),
	.full(fullProc75South),
	.dataIn(dataOutProc75South),
	.rd(rdProc88North),
	.empty(emptyProc88North),
	.dataOut(dataInProc88North));

	//FIFO 89 TO 88 
fifo fifo_proc89_to_proc88(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc89West),
	.full(fullProc89West),
	.dataIn(dataOutProc89West),
	.rd(rdProc88East),
	.empty(emptyProc88East),
	.dataOut(dataInProc88East));
	
	//FIFO 88 TO 89
fifo fifo_proc88_to_proc89(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc88East),
	.full(fullProc88East),
	.dataIn(dataOutProc88East),
	.rd(rdProc89West),
	.empty(emptyProc89West),
	.dataOut(dataInProc89West));
	
	//FIFO 89 TO 76 
fifo fifo_proc89_to_proc76(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc89North),
	.full(fullProc89North),
	.dataIn(dataOutProc89North),
	.rd(rdProc76South),
	.empty(emptyProc76South),
	.dataOut(dataInProc76South));
	
	//FIFO 76 TO 89
fifo fifo_proc76_to_proc89(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc76South),
	.full(fullProc76South),
	.dataIn(dataOutProc76South),
	.rd(rdProc89North),
	.empty(emptyProc89North),
	.dataOut(dataInProc89North));

	//FIFO 90 TO 89 
fifo fifo_proc90_to_proc89(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc90West),
	.full(fullProc90West),
	.dataIn(dataOutProc90West),
	.rd(rdProc89East),
	.empty(emptyProc89East),
	.dataOut(dataInProc89East));
	
	//FIFO 89 TO 90
fifo fifo_proc89_to_proc90(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc89East),
	.full(fullProc89East),
	.dataIn(dataOutProc89East),
	.rd(rdProc90West),
	.empty(emptyProc90West),
	.dataOut(dataInProc90West));
	
	//FIFO 90 TO 77 
fifo fifo_proc90_to_proc77(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc90North),
	.full(fullProc90North),
	.dataIn(dataOutProc90North),
	.rd(rdProc77South),
	.empty(emptyProc77South),
	.dataOut(dataInProc77South));
	
	//FIFO 77 TO 90
fifo fifo_proc77_to_proc90(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc77South),
	.full(fullProc77South),
	.dataIn(dataOutProc77South),
	.rd(rdProc90North),
	.empty(emptyProc90North),
	.dataOut(dataInProc90North));

	//FIFO 91 TO 78 
fifo fifo_proc91_to_proc78(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc91North),
	.full(fullProc91North),
	.dataIn(dataOutProc91North),
	.rd(rdProc78South),
	.empty(emptyProc78South),
	.dataOut(dataInProc78South));
	
	//FIFO 78 TO 91
fifo fifo_proc78_to_proc91(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc78South),
	.full(fullProc78South),
	.dataIn(dataOutProc78South),
	.rd(rdProc91North),
	.empty(emptyProc91North),
	.dataOut(dataInProc91North));

	//FIFO 92 TO 91 
fifo fifo_proc92_to_proc91(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc92West),
	.full(fullProc92West),
	.dataIn(dataOutProc92West),
	.rd(rdProc91East),
	.empty(emptyProc91East),
	.dataOut(dataInProc91East));
	
	//FIFO 91 TO 92
fifo fifo_proc91_to_proc92(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc91East),
	.full(fullProc91East),
	.dataIn(dataOutProc91East),
	.rd(rdProc92West),
	.empty(emptyProc92West),
	.dataOut(dataInProc92West));
	
	//FIFO 92 TO 79 
fifo fifo_proc92_to_proc79(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc92North),
	.full(fullProc92North),
	.dataIn(dataOutProc92North),
	.rd(rdProc79South),
	.empty(emptyProc79South),
	.dataOut(dataInProc79South));
	
	//FIFO 79 TO 92
fifo fifo_proc79_to_proc92(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc79South),
	.full(fullProc79South),
	.dataIn(dataOutProc79South),
	.rd(rdProc92North),
	.empty(emptyProc92North),
	.dataOut(dataInProc92North));

	//FIFO 93 TO 92 
fifo fifo_proc93_to_proc92(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc93West),
	.full(fullProc93West),
	.dataIn(dataOutProc93West),
	.rd(rdProc92East),
	.empty(emptyProc92East),
	.dataOut(dataInProc92East));
	
	//FIFO 92 TO 93
fifo fifo_proc92_to_proc93(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc92East),
	.full(fullProc92East),
	.dataIn(dataOutProc92East),
	.rd(rdProc93West),
	.empty(emptyProc93West),
	.dataOut(dataInProc93West));
	
	//FIFO 93 TO 80 
fifo fifo_proc93_to_proc80(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc93North),
	.full(fullProc93North),
	.dataIn(dataOutProc93North),
	.rd(rdProc80South),
	.empty(emptyProc80South),
	.dataOut(dataInProc80South));
	
	//FIFO 80 TO 93
fifo fifo_proc80_to_proc93(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc80South),
	.full(fullProc80South),
	.dataIn(dataOutProc80South),
	.rd(rdProc93North),
	.empty(emptyProc93North),
	.dataOut(dataInProc93North));

	//FIFO 94 TO 93 
fifo fifo_proc94_to_proc93(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc94West),
	.full(fullProc94West),
	.dataIn(dataOutProc94West),
	.rd(rdProc93East),
	.empty(emptyProc93East),
	.dataOut(dataInProc93East));
	
	//FIFO 93 TO 94
fifo fifo_proc93_to_proc94(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc93East),
	.full(fullProc93East),
	.dataIn(dataOutProc93East),
	.rd(rdProc94West),
	.empty(emptyProc94West),
	.dataOut(dataInProc94West));
	
	//FIFO 94 TO 81 
fifo fifo_proc94_to_proc81(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc94North),
	.full(fullProc94North),
	.dataIn(dataOutProc94North),
	.rd(rdProc81South),
	.empty(emptyProc81South),
	.dataOut(dataInProc81South));
	
	//FIFO 81 TO 94
fifo fifo_proc81_to_proc94(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc81South),
	.full(fullProc81South),
	.dataIn(dataOutProc81South),
	.rd(rdProc94North),
	.empty(emptyProc94North),
	.dataOut(dataInProc94North));

	//FIFO 95 TO 94 
fifo fifo_proc95_to_proc94(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc95West),
	.full(fullProc95West),
	.dataIn(dataOutProc95West),
	.rd(rdProc94East),
	.empty(emptyProc94East),
	.dataOut(dataInProc94East));
	
	//FIFO 94 TO 95
fifo fifo_proc94_to_proc95(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc94East),
	.full(fullProc94East),
	.dataIn(dataOutProc94East),
	.rd(rdProc95West),
	.empty(emptyProc95West),
	.dataOut(dataInProc95West));
	
	//FIFO 95 TO 82 
fifo fifo_proc95_to_proc82(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc95North),
	.full(fullProc95North),
	.dataIn(dataOutProc95North),
	.rd(rdProc82South),
	.empty(emptyProc82South),
	.dataOut(dataInProc82South));
	
	//FIFO 82 TO 95
fifo fifo_proc82_to_proc95(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc82South),
	.full(fullProc82South),
	.dataIn(dataOutProc82South),
	.rd(rdProc95North),
	.empty(emptyProc95North),
	.dataOut(dataInProc95North));

	//FIFO 96 TO 95 
fifo fifo_proc96_to_proc95(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc96West),
	.full(fullProc96West),
	.dataIn(dataOutProc96West),
	.rd(rdProc95East),
	.empty(emptyProc95East),
	.dataOut(dataInProc95East));
	
	//FIFO 95 TO 96
fifo fifo_proc95_to_proc96(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc95East),
	.full(fullProc95East),
	.dataIn(dataOutProc95East),
	.rd(rdProc96West),
	.empty(emptyProc96West),
	.dataOut(dataInProc96West));
	
	//FIFO 96 TO 83 
fifo fifo_proc96_to_proc83(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc96North),
	.full(fullProc96North),
	.dataIn(dataOutProc96North),
	.rd(rdProc83South),
	.empty(emptyProc83South),
	.dataOut(dataInProc83South));
	
	//FIFO 83 TO 96
fifo fifo_proc83_to_proc96(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc83South),
	.full(fullProc83South),
	.dataIn(dataOutProc83South),
	.rd(rdProc96North),
	.empty(emptyProc96North),
	.dataOut(dataInProc96North));

	//FIFO 97 TO 96 
fifo fifo_proc97_to_proc96(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc97West),
	.full(fullProc97West),
	.dataIn(dataOutProc97West),
	.rd(rdProc96East),
	.empty(emptyProc96East),
	.dataOut(dataInProc96East));
	
	//FIFO 96 TO 97
fifo fifo_proc96_to_proc97(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc96East),
	.full(fullProc96East),
	.dataIn(dataOutProc96East),
	.rd(rdProc97West),
	.empty(emptyProc97West),
	.dataOut(dataInProc97West));
	
	//FIFO 97 TO 84 
fifo fifo_proc97_to_proc84(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc97North),
	.full(fullProc97North),
	.dataIn(dataOutProc97North),
	.rd(rdProc84South),
	.empty(emptyProc84South),
	.dataOut(dataInProc84South));
	
	//FIFO 84 TO 97
fifo fifo_proc84_to_proc97(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc84South),
	.full(fullProc84South),
	.dataIn(dataOutProc84South),
	.rd(rdProc97North),
	.empty(emptyProc97North),
	.dataOut(dataInProc97North));

	//FIFO 98 TO 97 
fifo fifo_proc98_to_proc97(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc98West),
	.full(fullProc98West),
	.dataIn(dataOutProc98West),
	.rd(rdProc97East),
	.empty(emptyProc97East),
	.dataOut(dataInProc97East));
	
	//FIFO 97 TO 98
fifo fifo_proc97_to_proc98(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc97East),
	.full(fullProc97East),
	.dataIn(dataOutProc97East),
	.rd(rdProc98West),
	.empty(emptyProc98West),
	.dataOut(dataInProc98West));
	
	//FIFO 98 TO 85 
fifo fifo_proc98_to_proc85(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc98North),
	.full(fullProc98North),
	.dataIn(dataOutProc98North),
	.rd(rdProc85South),
	.empty(emptyProc85South),
	.dataOut(dataInProc85South));
	
	//FIFO 85 TO 98
fifo fifo_proc85_to_proc98(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc85South),
	.full(fullProc85South),
	.dataIn(dataOutProc85South),
	.rd(rdProc98North),
	.empty(emptyProc98North),
	.dataOut(dataInProc98North));

	//FIFO 99 TO 98 
fifo fifo_proc99_to_proc98(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc99West),
	.full(fullProc99West),
	.dataIn(dataOutProc99West),
	.rd(rdProc98East),
	.empty(emptyProc98East),
	.dataOut(dataInProc98East));
	
	//FIFO 98 TO 99
fifo fifo_proc98_to_proc99(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc98East),
	.full(fullProc98East),
	.dataIn(dataOutProc98East),
	.rd(rdProc99West),
	.empty(emptyProc99West),
	.dataOut(dataInProc99West));
	
	//FIFO 99 TO 86 
fifo fifo_proc99_to_proc86(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc99North),
	.full(fullProc99North),
	.dataIn(dataOutProc99North),
	.rd(rdProc86South),
	.empty(emptyProc86South),
	.dataOut(dataInProc86South));
	
	//FIFO 86 TO 99
fifo fifo_proc86_to_proc99(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc86South),
	.full(fullProc86South),
	.dataIn(dataOutProc86South),
	.rd(rdProc99North),
	.empty(emptyProc99North),
	.dataOut(dataInProc99North));

	//FIFO 100 TO 99 
fifo fifo_proc100_to_proc99(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc100West),
	.full(fullProc100West),
	.dataIn(dataOutProc100West),
	.rd(rdProc99East),
	.empty(emptyProc99East),
	.dataOut(dataInProc99East));
	
	//FIFO 99 TO 100
fifo fifo_proc99_to_proc100(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc99East),
	.full(fullProc99East),
	.dataIn(dataOutProc99East),
	.rd(rdProc100West),
	.empty(emptyProc100West),
	.dataOut(dataInProc100West));
	
	//FIFO 100 TO 87 
fifo fifo_proc100_to_proc87(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc100North),
	.full(fullProc100North),
	.dataIn(dataOutProc100North),
	.rd(rdProc87South),
	.empty(emptyProc87South),
	.dataOut(dataInProc87South));
	
	//FIFO 87 TO 100
fifo fifo_proc87_to_proc100(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc87South),
	.full(fullProc87South),
	.dataIn(dataOutProc87South),
	.rd(rdProc100North),
	.empty(emptyProc100North),
	.dataOut(dataInProc100North));

	//FIFO 101 TO 100 
fifo fifo_proc101_to_proc100(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc101West),
	.full(fullProc101West),
	.dataIn(dataOutProc101West),
	.rd(rdProc100East),
	.empty(emptyProc100East),
	.dataOut(dataInProc100East));
	
	//FIFO 100 TO 101
fifo fifo_proc100_to_proc101(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc100East),
	.full(fullProc100East),
	.dataIn(dataOutProc100East),
	.rd(rdProc101West),
	.empty(emptyProc101West),
	.dataOut(dataInProc101West));
	
	//FIFO 101 TO 88 
fifo fifo_proc101_to_proc88(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc101North),
	.full(fullProc101North),
	.dataIn(dataOutProc101North),
	.rd(rdProc88South),
	.empty(emptyProc88South),
	.dataOut(dataInProc88South));
	
	//FIFO 88 TO 101
fifo fifo_proc88_to_proc101(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc88South),
	.full(fullProc88South),
	.dataIn(dataOutProc88South),
	.rd(rdProc101North),
	.empty(emptyProc101North),
	.dataOut(dataInProc101North));

	//FIFO 102 TO 101 
fifo fifo_proc102_to_proc101(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc102West),
	.full(fullProc102West),
	.dataIn(dataOutProc102West),
	.rd(rdProc101East),
	.empty(emptyProc101East),
	.dataOut(dataInProc101East));
	
	//FIFO 101 TO 102
fifo fifo_proc101_to_proc102(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc101East),
	.full(fullProc101East),
	.dataIn(dataOutProc101East),
	.rd(rdProc102West),
	.empty(emptyProc102West),
	.dataOut(dataInProc102West));
	
	//FIFO 102 TO 89 
fifo fifo_proc102_to_proc89(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc102North),
	.full(fullProc102North),
	.dataIn(dataOutProc102North),
	.rd(rdProc89South),
	.empty(emptyProc89South),
	.dataOut(dataInProc89South));
	
	//FIFO 89 TO 102
fifo fifo_proc89_to_proc102(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc89South),
	.full(fullProc89South),
	.dataIn(dataOutProc89South),
	.rd(rdProc102North),
	.empty(emptyProc102North),
	.dataOut(dataInProc102North));

	//FIFO 103 TO 102 
fifo fifo_proc103_to_proc102(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc103West),
	.full(fullProc103West),
	.dataIn(dataOutProc103West),
	.rd(rdProc102East),
	.empty(emptyProc102East),
	.dataOut(dataInProc102East));
	
	//FIFO 102 TO 103
fifo fifo_proc102_to_proc103(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc102East),
	.full(fullProc102East),
	.dataIn(dataOutProc102East),
	.rd(rdProc103West),
	.empty(emptyProc103West),
	.dataOut(dataInProc103West));
	
	//FIFO 103 TO 90 
fifo fifo_proc103_to_proc90(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc103North),
	.full(fullProc103North),
	.dataIn(dataOutProc103North),
	.rd(rdProc90South),
	.empty(emptyProc90South),
	.dataOut(dataInProc90South));
	
	//FIFO 90 TO 103
fifo fifo_proc90_to_proc103(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc90South),
	.full(fullProc90South),
	.dataIn(dataOutProc90South),
	.rd(rdProc103North),
	.empty(emptyProc103North),
	.dataOut(dataInProc103North));

	//FIFO 104 TO 91 
fifo fifo_proc104_to_proc91(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc104North),
	.full(fullProc104North),
	.dataIn(dataOutProc104North),
	.rd(rdProc91South),
	.empty(emptyProc91South),
	.dataOut(dataInProc91South));
	
	//FIFO 91 TO 104
fifo fifo_proc91_to_proc104(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc91South),
	.full(fullProc91South),
	.dataIn(dataOutProc91South),
	.rd(rdProc104North),
	.empty(emptyProc104North),
	.dataOut(dataInProc104North));

	//FIFO 105 TO 104 
fifo fifo_proc105_to_proc104(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc105West),
	.full(fullProc105West),
	.dataIn(dataOutProc105West),
	.rd(rdProc104East),
	.empty(emptyProc104East),
	.dataOut(dataInProc104East));
	
	//FIFO 104 TO 105
fifo fifo_proc104_to_proc105(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc104East),
	.full(fullProc104East),
	.dataIn(dataOutProc104East),
	.rd(rdProc105West),
	.empty(emptyProc105West),
	.dataOut(dataInProc105West));
	
	//FIFO 105 TO 92 
fifo fifo_proc105_to_proc92(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc105North),
	.full(fullProc105North),
	.dataIn(dataOutProc105North),
	.rd(rdProc92South),
	.empty(emptyProc92South),
	.dataOut(dataInProc92South));
	
	//FIFO 92 TO 105
fifo fifo_proc92_to_proc105(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc92South),
	.full(fullProc92South),
	.dataIn(dataOutProc92South),
	.rd(rdProc105North),
	.empty(emptyProc105North),
	.dataOut(dataInProc105North));

	//FIFO 106 TO 105 
fifo fifo_proc106_to_proc105(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc106West),
	.full(fullProc106West),
	.dataIn(dataOutProc106West),
	.rd(rdProc105East),
	.empty(emptyProc105East),
	.dataOut(dataInProc105East));
	
	//FIFO 105 TO 106
fifo fifo_proc105_to_proc106(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc105East),
	.full(fullProc105East),
	.dataIn(dataOutProc105East),
	.rd(rdProc106West),
	.empty(emptyProc106West),
	.dataOut(dataInProc106West));
	
	//FIFO 106 TO 93 
fifo fifo_proc106_to_proc93(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc106North),
	.full(fullProc106North),
	.dataIn(dataOutProc106North),
	.rd(rdProc93South),
	.empty(emptyProc93South),
	.dataOut(dataInProc93South));
	
	//FIFO 93 TO 106
fifo fifo_proc93_to_proc106(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc93South),
	.full(fullProc93South),
	.dataIn(dataOutProc93South),
	.rd(rdProc106North),
	.empty(emptyProc106North),
	.dataOut(dataInProc106North));

	//FIFO 107 TO 106 
fifo fifo_proc107_to_proc106(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc107West),
	.full(fullProc107West),
	.dataIn(dataOutProc107West),
	.rd(rdProc106East),
	.empty(emptyProc106East),
	.dataOut(dataInProc106East));
	
	//FIFO 106 TO 107
fifo fifo_proc106_to_proc107(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc106East),
	.full(fullProc106East),
	.dataIn(dataOutProc106East),
	.rd(rdProc107West),
	.empty(emptyProc107West),
	.dataOut(dataInProc107West));
	
	//FIFO 107 TO 94 
fifo fifo_proc107_to_proc94(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc107North),
	.full(fullProc107North),
	.dataIn(dataOutProc107North),
	.rd(rdProc94South),
	.empty(emptyProc94South),
	.dataOut(dataInProc94South));
	
	//FIFO 94 TO 107
fifo fifo_proc94_to_proc107(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc94South),
	.full(fullProc94South),
	.dataIn(dataOutProc94South),
	.rd(rdProc107North),
	.empty(emptyProc107North),
	.dataOut(dataInProc107North));

	//FIFO 108 TO 107 
fifo fifo_proc108_to_proc107(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc108West),
	.full(fullProc108West),
	.dataIn(dataOutProc108West),
	.rd(rdProc107East),
	.empty(emptyProc107East),
	.dataOut(dataInProc107East));
	
	//FIFO 107 TO 108
fifo fifo_proc107_to_proc108(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc107East),
	.full(fullProc107East),
	.dataIn(dataOutProc107East),
	.rd(rdProc108West),
	.empty(emptyProc108West),
	.dataOut(dataInProc108West));
	
	//FIFO 108 TO 95 
fifo fifo_proc108_to_proc95(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc108North),
	.full(fullProc108North),
	.dataIn(dataOutProc108North),
	.rd(rdProc95South),
	.empty(emptyProc95South),
	.dataOut(dataInProc95South));
	
	//FIFO 95 TO 108
fifo fifo_proc95_to_proc108(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc95South),
	.full(fullProc95South),
	.dataIn(dataOutProc95South),
	.rd(rdProc108North),
	.empty(emptyProc108North),
	.dataOut(dataInProc108North));

	//FIFO 109 TO 108 
fifo fifo_proc109_to_proc108(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc109West),
	.full(fullProc109West),
	.dataIn(dataOutProc109West),
	.rd(rdProc108East),
	.empty(emptyProc108East),
	.dataOut(dataInProc108East));
	
	//FIFO 108 TO 109
fifo fifo_proc108_to_proc109(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc108East),
	.full(fullProc108East),
	.dataIn(dataOutProc108East),
	.rd(rdProc109West),
	.empty(emptyProc109West),
	.dataOut(dataInProc109West));
	
	//FIFO 109 TO 96 
fifo fifo_proc109_to_proc96(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc109North),
	.full(fullProc109North),
	.dataIn(dataOutProc109North),
	.rd(rdProc96South),
	.empty(emptyProc96South),
	.dataOut(dataInProc96South));
	
	//FIFO 96 TO 109
fifo fifo_proc96_to_proc109(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc96South),
	.full(fullProc96South),
	.dataIn(dataOutProc96South),
	.rd(rdProc109North),
	.empty(emptyProc109North),
	.dataOut(dataInProc109North));

	//FIFO 110 TO 109 
fifo fifo_proc110_to_proc109(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc110West),
	.full(fullProc110West),
	.dataIn(dataOutProc110West),
	.rd(rdProc109East),
	.empty(emptyProc109East),
	.dataOut(dataInProc109East));
	
	//FIFO 109 TO 110
fifo fifo_proc109_to_proc110(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc109East),
	.full(fullProc109East),
	.dataIn(dataOutProc109East),
	.rd(rdProc110West),
	.empty(emptyProc110West),
	.dataOut(dataInProc110West));
	
	//FIFO 110 TO 97 
fifo fifo_proc110_to_proc97(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc110North),
	.full(fullProc110North),
	.dataIn(dataOutProc110North),
	.rd(rdProc97South),
	.empty(emptyProc97South),
	.dataOut(dataInProc97South));
	
	//FIFO 97 TO 110
fifo fifo_proc97_to_proc110(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc97South),
	.full(fullProc97South),
	.dataIn(dataOutProc97South),
	.rd(rdProc110North),
	.empty(emptyProc110North),
	.dataOut(dataInProc110North));

	//FIFO 111 TO 110 
fifo fifo_proc111_to_proc110(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc111West),
	.full(fullProc111West),
	.dataIn(dataOutProc111West),
	.rd(rdProc110East),
	.empty(emptyProc110East),
	.dataOut(dataInProc110East));
	
	//FIFO 110 TO 111
fifo fifo_proc110_to_proc111(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc110East),
	.full(fullProc110East),
	.dataIn(dataOutProc110East),
	.rd(rdProc111West),
	.empty(emptyProc111West),
	.dataOut(dataInProc111West));
	
	//FIFO 111 TO 98 
fifo fifo_proc111_to_proc98(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc111North),
	.full(fullProc111North),
	.dataIn(dataOutProc111North),
	.rd(rdProc98South),
	.empty(emptyProc98South),
	.dataOut(dataInProc98South));
	
	//FIFO 98 TO 111
fifo fifo_proc98_to_proc111(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc98South),
	.full(fullProc98South),
	.dataIn(dataOutProc98South),
	.rd(rdProc111North),
	.empty(emptyProc111North),
	.dataOut(dataInProc111North));

	//FIFO 112 TO 111 
fifo fifo_proc112_to_proc111(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc112West),
	.full(fullProc112West),
	.dataIn(dataOutProc112West),
	.rd(rdProc111East),
	.empty(emptyProc111East),
	.dataOut(dataInProc111East));
	
	//FIFO 111 TO 112
fifo fifo_proc111_to_proc112(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc111East),
	.full(fullProc111East),
	.dataIn(dataOutProc111East),
	.rd(rdProc112West),
	.empty(emptyProc112West),
	.dataOut(dataInProc112West));
	
	//FIFO 112 TO 99 
fifo fifo_proc112_to_proc99(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc112North),
	.full(fullProc112North),
	.dataIn(dataOutProc112North),
	.rd(rdProc99South),
	.empty(emptyProc99South),
	.dataOut(dataInProc99South));
	
	//FIFO 99 TO 112
fifo fifo_proc99_to_proc112(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc99South),
	.full(fullProc99South),
	.dataIn(dataOutProc99South),
	.rd(rdProc112North),
	.empty(emptyProc112North),
	.dataOut(dataInProc112North));

	//FIFO 113 TO 112 
fifo fifo_proc113_to_proc112(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc113West),
	.full(fullProc113West),
	.dataIn(dataOutProc113West),
	.rd(rdProc112East),
	.empty(emptyProc112East),
	.dataOut(dataInProc112East));
	
	//FIFO 112 TO 113
fifo fifo_proc112_to_proc113(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc112East),
	.full(fullProc112East),
	.dataIn(dataOutProc112East),
	.rd(rdProc113West),
	.empty(emptyProc113West),
	.dataOut(dataInProc113West));
	
	//FIFO 113 TO 100 
fifo fifo_proc113_to_proc100(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc113North),
	.full(fullProc113North),
	.dataIn(dataOutProc113North),
	.rd(rdProc100South),
	.empty(emptyProc100South),
	.dataOut(dataInProc100South));
	
	//FIFO 100 TO 113
fifo fifo_proc100_to_proc113(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc100South),
	.full(fullProc100South),
	.dataIn(dataOutProc100South),
	.rd(rdProc113North),
	.empty(emptyProc113North),
	.dataOut(dataInProc113North));

	//FIFO 114 TO 113 
fifo fifo_proc114_to_proc113(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc114West),
	.full(fullProc114West),
	.dataIn(dataOutProc114West),
	.rd(rdProc113East),
	.empty(emptyProc113East),
	.dataOut(dataInProc113East));
	
	//FIFO 113 TO 114
fifo fifo_proc113_to_proc114(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc113East),
	.full(fullProc113East),
	.dataIn(dataOutProc113East),
	.rd(rdProc114West),
	.empty(emptyProc114West),
	.dataOut(dataInProc114West));
	
	//FIFO 114 TO 101 
fifo fifo_proc114_to_proc101(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc114North),
	.full(fullProc114North),
	.dataIn(dataOutProc114North),
	.rd(rdProc101South),
	.empty(emptyProc101South),
	.dataOut(dataInProc101South));
	
	//FIFO 101 TO 114
fifo fifo_proc101_to_proc114(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc101South),
	.full(fullProc101South),
	.dataIn(dataOutProc101South),
	.rd(rdProc114North),
	.empty(emptyProc114North),
	.dataOut(dataInProc114North));

	//FIFO 115 TO 114 
fifo fifo_proc115_to_proc114(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc115West),
	.full(fullProc115West),
	.dataIn(dataOutProc115West),
	.rd(rdProc114East),
	.empty(emptyProc114East),
	.dataOut(dataInProc114East));
	
	//FIFO 114 TO 115
fifo fifo_proc114_to_proc115(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc114East),
	.full(fullProc114East),
	.dataIn(dataOutProc114East),
	.rd(rdProc115West),
	.empty(emptyProc115West),
	.dataOut(dataInProc115West));
	
	//FIFO 115 TO 102 
fifo fifo_proc115_to_proc102(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc115North),
	.full(fullProc115North),
	.dataIn(dataOutProc115North),
	.rd(rdProc102South),
	.empty(emptyProc102South),
	.dataOut(dataInProc102South));
	
	//FIFO 102 TO 115
fifo fifo_proc102_to_proc115(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc102South),
	.full(fullProc102South),
	.dataIn(dataOutProc102South),
	.rd(rdProc115North),
	.empty(emptyProc115North),
	.dataOut(dataInProc115North));

	//FIFO 116 TO 115 
fifo fifo_proc116_to_proc115(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc116West),
	.full(fullProc116West),
	.dataIn(dataOutProc116West),
	.rd(rdProc115East),
	.empty(emptyProc115East),
	.dataOut(dataInProc115East));
	
	//FIFO 115 TO 116
fifo fifo_proc115_to_proc116(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc115East),
	.full(fullProc115East),
	.dataIn(dataOutProc115East),
	.rd(rdProc116West),
	.empty(emptyProc116West),
	.dataOut(dataInProc116West));
	
	//FIFO 116 TO 103 
fifo fifo_proc116_to_proc103(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc116North),
	.full(fullProc116North),
	.dataIn(dataOutProc116North),
	.rd(rdProc103South),
	.empty(emptyProc103South),
	.dataOut(dataInProc103South));
	
	//FIFO 103 TO 116
fifo fifo_proc103_to_proc116(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc103South),
	.full(fullProc103South),
	.dataIn(dataOutProc103South),
	.rd(rdProc116North),
	.empty(emptyProc116North),
	.dataOut(dataInProc116North));

	//FIFO 117 TO 104 
fifo fifo_proc117_to_proc104(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc117North),
	.full(fullProc117North),
	.dataIn(dataOutProc117North),
	.rd(rdProc104South),
	.empty(emptyProc104South),
	.dataOut(dataInProc104South));
	
	//FIFO 104 TO 117
fifo fifo_proc104_to_proc117(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc104South),
	.full(fullProc104South),
	.dataIn(dataOutProc104South),
	.rd(rdProc117North),
	.empty(emptyProc117North),
	.dataOut(dataInProc117North));

	//FIFO 118 TO 117 
fifo fifo_proc118_to_proc117(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc118West),
	.full(fullProc118West),
	.dataIn(dataOutProc118West),
	.rd(rdProc117East),
	.empty(emptyProc117East),
	.dataOut(dataInProc117East));
	
	//FIFO 117 TO 118
fifo fifo_proc117_to_proc118(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc117East),
	.full(fullProc117East),
	.dataIn(dataOutProc117East),
	.rd(rdProc118West),
	.empty(emptyProc118West),
	.dataOut(dataInProc118West));
	
	//FIFO 118 TO 105 
fifo fifo_proc118_to_proc105(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc118North),
	.full(fullProc118North),
	.dataIn(dataOutProc118North),
	.rd(rdProc105South),
	.empty(emptyProc105South),
	.dataOut(dataInProc105South));
	
	//FIFO 105 TO 118
fifo fifo_proc105_to_proc118(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc105South),
	.full(fullProc105South),
	.dataIn(dataOutProc105South),
	.rd(rdProc118North),
	.empty(emptyProc118North),
	.dataOut(dataInProc118North));

	//FIFO 119 TO 118 
fifo fifo_proc119_to_proc118(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc119West),
	.full(fullProc119West),
	.dataIn(dataOutProc119West),
	.rd(rdProc118East),
	.empty(emptyProc118East),
	.dataOut(dataInProc118East));
	
	//FIFO 118 TO 119
fifo fifo_proc118_to_proc119(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc118East),
	.full(fullProc118East),
	.dataIn(dataOutProc118East),
	.rd(rdProc119West),
	.empty(emptyProc119West),
	.dataOut(dataInProc119West));
	
	//FIFO 119 TO 106 
fifo fifo_proc119_to_proc106(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc119North),
	.full(fullProc119North),
	.dataIn(dataOutProc119North),
	.rd(rdProc106South),
	.empty(emptyProc106South),
	.dataOut(dataInProc106South));
	
	//FIFO 106 TO 119
fifo fifo_proc106_to_proc119(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc106South),
	.full(fullProc106South),
	.dataIn(dataOutProc106South),
	.rd(rdProc119North),
	.empty(emptyProc119North),
	.dataOut(dataInProc119North));

	//FIFO 120 TO 119 
fifo fifo_proc120_to_proc119(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc120West),
	.full(fullProc120West),
	.dataIn(dataOutProc120West),
	.rd(rdProc119East),
	.empty(emptyProc119East),
	.dataOut(dataInProc119East));
	
	//FIFO 119 TO 120
fifo fifo_proc119_to_proc120(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc119East),
	.full(fullProc119East),
	.dataIn(dataOutProc119East),
	.rd(rdProc120West),
	.empty(emptyProc120West),
	.dataOut(dataInProc120West));
	
	//FIFO 120 TO 107 
fifo fifo_proc120_to_proc107(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc120North),
	.full(fullProc120North),
	.dataIn(dataOutProc120North),
	.rd(rdProc107South),
	.empty(emptyProc107South),
	.dataOut(dataInProc107South));
	
	//FIFO 107 TO 120
fifo fifo_proc107_to_proc120(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc107South),
	.full(fullProc107South),
	.dataIn(dataOutProc107South),
	.rd(rdProc120North),
	.empty(emptyProc120North),
	.dataOut(dataInProc120North));

	//FIFO 121 TO 120 
fifo fifo_proc121_to_proc120(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc121West),
	.full(fullProc121West),
	.dataIn(dataOutProc121West),
	.rd(rdProc120East),
	.empty(emptyProc120East),
	.dataOut(dataInProc120East));
	
	//FIFO 120 TO 121
fifo fifo_proc120_to_proc121(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc120East),
	.full(fullProc120East),
	.dataIn(dataOutProc120East),
	.rd(rdProc121West),
	.empty(emptyProc121West),
	.dataOut(dataInProc121West));
	
	//FIFO 121 TO 108 
fifo fifo_proc121_to_proc108(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc121North),
	.full(fullProc121North),
	.dataIn(dataOutProc121North),
	.rd(rdProc108South),
	.empty(emptyProc108South),
	.dataOut(dataInProc108South));
	
	//FIFO 108 TO 121
fifo fifo_proc108_to_proc121(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc108South),
	.full(fullProc108South),
	.dataIn(dataOutProc108South),
	.rd(rdProc121North),
	.empty(emptyProc121North),
	.dataOut(dataInProc121North));

	//FIFO 122 TO 121 
fifo fifo_proc122_to_proc121(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc122West),
	.full(fullProc122West),
	.dataIn(dataOutProc122West),
	.rd(rdProc121East),
	.empty(emptyProc121East),
	.dataOut(dataInProc121East));
	
	//FIFO 121 TO 122
fifo fifo_proc121_to_proc122(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc121East),
	.full(fullProc121East),
	.dataIn(dataOutProc121East),
	.rd(rdProc122West),
	.empty(emptyProc122West),
	.dataOut(dataInProc122West));
	
	//FIFO 122 TO 109 
fifo fifo_proc122_to_proc109(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc122North),
	.full(fullProc122North),
	.dataIn(dataOutProc122North),
	.rd(rdProc109South),
	.empty(emptyProc109South),
	.dataOut(dataInProc109South));
	
	//FIFO 109 TO 122
fifo fifo_proc109_to_proc122(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc109South),
	.full(fullProc109South),
	.dataIn(dataOutProc109South),
	.rd(rdProc122North),
	.empty(emptyProc122North),
	.dataOut(dataInProc122North));

	//FIFO 123 TO 122 
fifo fifo_proc123_to_proc122(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc123West),
	.full(fullProc123West),
	.dataIn(dataOutProc123West),
	.rd(rdProc122East),
	.empty(emptyProc122East),
	.dataOut(dataInProc122East));
	
	//FIFO 122 TO 123
fifo fifo_proc122_to_proc123(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc122East),
	.full(fullProc122East),
	.dataIn(dataOutProc122East),
	.rd(rdProc123West),
	.empty(emptyProc123West),
	.dataOut(dataInProc123West));
	
	//FIFO 123 TO 110 
fifo fifo_proc123_to_proc110(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc123North),
	.full(fullProc123North),
	.dataIn(dataOutProc123North),
	.rd(rdProc110South),
	.empty(emptyProc110South),
	.dataOut(dataInProc110South));
	
	//FIFO 110 TO 123
fifo fifo_proc110_to_proc123(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc110South),
	.full(fullProc110South),
	.dataIn(dataOutProc110South),
	.rd(rdProc123North),
	.empty(emptyProc123North),
	.dataOut(dataInProc123North));

	//FIFO 124 TO 123 
fifo fifo_proc124_to_proc123(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc124West),
	.full(fullProc124West),
	.dataIn(dataOutProc124West),
	.rd(rdProc123East),
	.empty(emptyProc123East),
	.dataOut(dataInProc123East));
	
	//FIFO 123 TO 124
fifo fifo_proc123_to_proc124(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc123East),
	.full(fullProc123East),
	.dataIn(dataOutProc123East),
	.rd(rdProc124West),
	.empty(emptyProc124West),
	.dataOut(dataInProc124West));
	
	//FIFO 124 TO 111 
fifo fifo_proc124_to_proc111(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc124North),
	.full(fullProc124North),
	.dataIn(dataOutProc124North),
	.rd(rdProc111South),
	.empty(emptyProc111South),
	.dataOut(dataInProc111South));
	
	//FIFO 111 TO 124
fifo fifo_proc111_to_proc124(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc111South),
	.full(fullProc111South),
	.dataIn(dataOutProc111South),
	.rd(rdProc124North),
	.empty(emptyProc124North),
	.dataOut(dataInProc124North));

	//FIFO 125 TO 124 
fifo fifo_proc125_to_proc124(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc125West),
	.full(fullProc125West),
	.dataIn(dataOutProc125West),
	.rd(rdProc124East),
	.empty(emptyProc124East),
	.dataOut(dataInProc124East));
	
	//FIFO 124 TO 125
fifo fifo_proc124_to_proc125(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc124East),
	.full(fullProc124East),
	.dataIn(dataOutProc124East),
	.rd(rdProc125West),
	.empty(emptyProc125West),
	.dataOut(dataInProc125West));
	
	//FIFO 125 TO 112 
fifo fifo_proc125_to_proc112(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc125North),
	.full(fullProc125North),
	.dataIn(dataOutProc125North),
	.rd(rdProc112South),
	.empty(emptyProc112South),
	.dataOut(dataInProc112South));
	
	//FIFO 112 TO 125
fifo fifo_proc112_to_proc125(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc112South),
	.full(fullProc112South),
	.dataIn(dataOutProc112South),
	.rd(rdProc125North),
	.empty(emptyProc125North),
	.dataOut(dataInProc125North));

	//FIFO 126 TO 125 
fifo fifo_proc126_to_proc125(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc126West),
	.full(fullProc126West),
	.dataIn(dataOutProc126West),
	.rd(rdProc125East),
	.empty(emptyProc125East),
	.dataOut(dataInProc125East));
	
	//FIFO 125 TO 126
fifo fifo_proc125_to_proc126(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc125East),
	.full(fullProc125East),
	.dataIn(dataOutProc125East),
	.rd(rdProc126West),
	.empty(emptyProc126West),
	.dataOut(dataInProc126West));
	
	//FIFO 126 TO 113 
fifo fifo_proc126_to_proc113(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc126North),
	.full(fullProc126North),
	.dataIn(dataOutProc126North),
	.rd(rdProc113South),
	.empty(emptyProc113South),
	.dataOut(dataInProc113South));
	
	//FIFO 113 TO 126
fifo fifo_proc113_to_proc126(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc113South),
	.full(fullProc113South),
	.dataIn(dataOutProc113South),
	.rd(rdProc126North),
	.empty(emptyProc126North),
	.dataOut(dataInProc126North));

	//FIFO 127 TO 126 
fifo fifo_proc127_to_proc126(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc127West),
	.full(fullProc127West),
	.dataIn(dataOutProc127West),
	.rd(rdProc126East),
	.empty(emptyProc126East),
	.dataOut(dataInProc126East));
	
	//FIFO 126 TO 127
fifo fifo_proc126_to_proc127(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc126East),
	.full(fullProc126East),
	.dataIn(dataOutProc126East),
	.rd(rdProc127West),
	.empty(emptyProc127West),
	.dataOut(dataInProc127West));
	
	//FIFO 127 TO 114 
fifo fifo_proc127_to_proc114(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc127North),
	.full(fullProc127North),
	.dataIn(dataOutProc127North),
	.rd(rdProc114South),
	.empty(emptyProc114South),
	.dataOut(dataInProc114South));
	
	//FIFO 114 TO 127
fifo fifo_proc114_to_proc127(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc114South),
	.full(fullProc114South),
	.dataIn(dataOutProc114South),
	.rd(rdProc127North),
	.empty(emptyProc127North),
	.dataOut(dataInProc127North));

	//FIFO 128 TO 127 
fifo fifo_proc128_to_proc127(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc128West),
	.full(fullProc128West),
	.dataIn(dataOutProc128West),
	.rd(rdProc127East),
	.empty(emptyProc127East),
	.dataOut(dataInProc127East));
	
	//FIFO 127 TO 128
fifo fifo_proc127_to_proc128(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc127East),
	.full(fullProc127East),
	.dataIn(dataOutProc127East),
	.rd(rdProc128West),
	.empty(emptyProc128West),
	.dataOut(dataInProc128West));
	
	//FIFO 128 TO 115 
fifo fifo_proc128_to_proc115(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc128North),
	.full(fullProc128North),
	.dataIn(dataOutProc128North),
	.rd(rdProc115South),
	.empty(emptyProc115South),
	.dataOut(dataInProc115South));
	
	//FIFO 115 TO 128
fifo fifo_proc115_to_proc128(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc115South),
	.full(fullProc115South),
	.dataIn(dataOutProc115South),
	.rd(rdProc128North),
	.empty(emptyProc128North),
	.dataOut(dataInProc128North));

	//FIFO 129 TO 128 
fifo fifo_proc129_to_proc128(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc129West),
	.full(fullProc129West),
	.dataIn(dataOutProc129West),
	.rd(rdProc128East),
	.empty(emptyProc128East),
	.dataOut(dataInProc128East));
	
	//FIFO 128 TO 129
fifo fifo_proc128_to_proc129(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc128East),
	.full(fullProc128East),
	.dataIn(dataOutProc128East),
	.rd(rdProc129West),
	.empty(emptyProc129West),
	.dataOut(dataInProc129West));
	
	//FIFO 129 TO 116 
fifo fifo_proc129_to_proc116(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc129North),
	.full(fullProc129North),
	.dataIn(dataOutProc129North),
	.rd(rdProc116South),
	.empty(emptyProc116South),
	.dataOut(dataInProc116South));
	
	//FIFO 116 TO 129
fifo fifo_proc116_to_proc129(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc116South),
	.full(fullProc116South),
	.dataIn(dataOutProc116South),
	.rd(rdProc129North),
	.empty(emptyProc129North),
	.dataOut(dataInProc129North));

	//FIFO 130 TO 117 
fifo fifo_proc130_to_proc117(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc130North),
	.full(fullProc130North),
	.dataIn(dataOutProc130North),
	.rd(rdProc117South),
	.empty(emptyProc117South),
	.dataOut(dataInProc117South));
	
	//FIFO 117 TO 130
fifo fifo_proc117_to_proc130(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc117South),
	.full(fullProc117South),
	.dataIn(dataOutProc117South),
	.rd(rdProc130North),
	.empty(emptyProc130North),
	.dataOut(dataInProc130North));

	//FIFO 131 TO 130 
fifo fifo_proc131_to_proc130(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc131West),
	.full(fullProc131West),
	.dataIn(dataOutProc131West),
	.rd(rdProc130East),
	.empty(emptyProc130East),
	.dataOut(dataInProc130East));
	
	//FIFO 130 TO 131
fifo fifo_proc130_to_proc131(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc130East),
	.full(fullProc130East),
	.dataIn(dataOutProc130East),
	.rd(rdProc131West),
	.empty(emptyProc131West),
	.dataOut(dataInProc131West));
	
	//FIFO 131 TO 118 
fifo fifo_proc131_to_proc118(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc131North),
	.full(fullProc131North),
	.dataIn(dataOutProc131North),
	.rd(rdProc118South),
	.empty(emptyProc118South),
	.dataOut(dataInProc118South));
	
	//FIFO 118 TO 131
fifo fifo_proc118_to_proc131(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc118South),
	.full(fullProc118South),
	.dataIn(dataOutProc118South),
	.rd(rdProc131North),
	.empty(emptyProc131North),
	.dataOut(dataInProc131North));

	//FIFO 132 TO 131 
fifo fifo_proc132_to_proc131(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc132West),
	.full(fullProc132West),
	.dataIn(dataOutProc132West),
	.rd(rdProc131East),
	.empty(emptyProc131East),
	.dataOut(dataInProc131East));
	
	//FIFO 131 TO 132
fifo fifo_proc131_to_proc132(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc131East),
	.full(fullProc131East),
	.dataIn(dataOutProc131East),
	.rd(rdProc132West),
	.empty(emptyProc132West),
	.dataOut(dataInProc132West));
	
	//FIFO 132 TO 119 
fifo fifo_proc132_to_proc119(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc132North),
	.full(fullProc132North),
	.dataIn(dataOutProc132North),
	.rd(rdProc119South),
	.empty(emptyProc119South),
	.dataOut(dataInProc119South));
	
	//FIFO 119 TO 132
fifo fifo_proc119_to_proc132(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc119South),
	.full(fullProc119South),
	.dataIn(dataOutProc119South),
	.rd(rdProc132North),
	.empty(emptyProc132North),
	.dataOut(dataInProc132North));

	//FIFO 133 TO 132 
fifo fifo_proc133_to_proc132(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc133West),
	.full(fullProc133West),
	.dataIn(dataOutProc133West),
	.rd(rdProc132East),
	.empty(emptyProc132East),
	.dataOut(dataInProc132East));
	
	//FIFO 132 TO 133
fifo fifo_proc132_to_proc133(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc132East),
	.full(fullProc132East),
	.dataIn(dataOutProc132East),
	.rd(rdProc133West),
	.empty(emptyProc133West),
	.dataOut(dataInProc133West));
	
	//FIFO 133 TO 120 
fifo fifo_proc133_to_proc120(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc133North),
	.full(fullProc133North),
	.dataIn(dataOutProc133North),
	.rd(rdProc120South),
	.empty(emptyProc120South),
	.dataOut(dataInProc120South));
	
	//FIFO 120 TO 133
fifo fifo_proc120_to_proc133(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc120South),
	.full(fullProc120South),
	.dataIn(dataOutProc120South),
	.rd(rdProc133North),
	.empty(emptyProc133North),
	.dataOut(dataInProc133North));

	//FIFO 134 TO 133 
fifo fifo_proc134_to_proc133(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc134West),
	.full(fullProc134West),
	.dataIn(dataOutProc134West),
	.rd(rdProc133East),
	.empty(emptyProc133East),
	.dataOut(dataInProc133East));
	
	//FIFO 133 TO 134
fifo fifo_proc133_to_proc134(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc133East),
	.full(fullProc133East),
	.dataIn(dataOutProc133East),
	.rd(rdProc134West),
	.empty(emptyProc134West),
	.dataOut(dataInProc134West));
	
	//FIFO 134 TO 121 
fifo fifo_proc134_to_proc121(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc134North),
	.full(fullProc134North),
	.dataIn(dataOutProc134North),
	.rd(rdProc121South),
	.empty(emptyProc121South),
	.dataOut(dataInProc121South));
	
	//FIFO 121 TO 134
fifo fifo_proc121_to_proc134(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc121South),
	.full(fullProc121South),
	.dataIn(dataOutProc121South),
	.rd(rdProc134North),
	.empty(emptyProc134North),
	.dataOut(dataInProc134North));

	//FIFO 135 TO 134 
fifo fifo_proc135_to_proc134(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc135West),
	.full(fullProc135West),
	.dataIn(dataOutProc135West),
	.rd(rdProc134East),
	.empty(emptyProc134East),
	.dataOut(dataInProc134East));
	
	//FIFO 134 TO 135
fifo fifo_proc134_to_proc135(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc134East),
	.full(fullProc134East),
	.dataIn(dataOutProc134East),
	.rd(rdProc135West),
	.empty(emptyProc135West),
	.dataOut(dataInProc135West));
	
	//FIFO 135 TO 122 
fifo fifo_proc135_to_proc122(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc135North),
	.full(fullProc135North),
	.dataIn(dataOutProc135North),
	.rd(rdProc122South),
	.empty(emptyProc122South),
	.dataOut(dataInProc122South));
	
	//FIFO 122 TO 135
fifo fifo_proc122_to_proc135(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc122South),
	.full(fullProc122South),
	.dataIn(dataOutProc122South),
	.rd(rdProc135North),
	.empty(emptyProc135North),
	.dataOut(dataInProc135North));

	//FIFO 136 TO 135 
fifo fifo_proc136_to_proc135(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc136West),
	.full(fullProc136West),
	.dataIn(dataOutProc136West),
	.rd(rdProc135East),
	.empty(emptyProc135East),
	.dataOut(dataInProc135East));
	
	//FIFO 135 TO 136
fifo fifo_proc135_to_proc136(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc135East),
	.full(fullProc135East),
	.dataIn(dataOutProc135East),
	.rd(rdProc136West),
	.empty(emptyProc136West),
	.dataOut(dataInProc136West));
	
	//FIFO 136 TO 123 
fifo fifo_proc136_to_proc123(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc136North),
	.full(fullProc136North),
	.dataIn(dataOutProc136North),
	.rd(rdProc123South),
	.empty(emptyProc123South),
	.dataOut(dataInProc123South));
	
	//FIFO 123 TO 136
fifo fifo_proc123_to_proc136(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc123South),
	.full(fullProc123South),
	.dataIn(dataOutProc123South),
	.rd(rdProc136North),
	.empty(emptyProc136North),
	.dataOut(dataInProc136North));

	//FIFO 137 TO 136 
fifo fifo_proc137_to_proc136(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc137West),
	.full(fullProc137West),
	.dataIn(dataOutProc137West),
	.rd(rdProc136East),
	.empty(emptyProc136East),
	.dataOut(dataInProc136East));
	
	//FIFO 136 TO 137
fifo fifo_proc136_to_proc137(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc136East),
	.full(fullProc136East),
	.dataIn(dataOutProc136East),
	.rd(rdProc137West),
	.empty(emptyProc137West),
	.dataOut(dataInProc137West));
	
	//FIFO 137 TO 124 
fifo fifo_proc137_to_proc124(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc137North),
	.full(fullProc137North),
	.dataIn(dataOutProc137North),
	.rd(rdProc124South),
	.empty(emptyProc124South),
	.dataOut(dataInProc124South));
	
	//FIFO 124 TO 137
fifo fifo_proc124_to_proc137(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc124South),
	.full(fullProc124South),
	.dataIn(dataOutProc124South),
	.rd(rdProc137North),
	.empty(emptyProc137North),
	.dataOut(dataInProc137North));

	//FIFO 138 TO 137 
fifo fifo_proc138_to_proc137(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc138West),
	.full(fullProc138West),
	.dataIn(dataOutProc138West),
	.rd(rdProc137East),
	.empty(emptyProc137East),
	.dataOut(dataInProc137East));
	
	//FIFO 137 TO 138
fifo fifo_proc137_to_proc138(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc137East),
	.full(fullProc137East),
	.dataIn(dataOutProc137East),
	.rd(rdProc138West),
	.empty(emptyProc138West),
	.dataOut(dataInProc138West));
	
	//FIFO 138 TO 125 
fifo fifo_proc138_to_proc125(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc138North),
	.full(fullProc138North),
	.dataIn(dataOutProc138North),
	.rd(rdProc125South),
	.empty(emptyProc125South),
	.dataOut(dataInProc125South));
	
	//FIFO 125 TO 138
fifo fifo_proc125_to_proc138(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc125South),
	.full(fullProc125South),
	.dataIn(dataOutProc125South),
	.rd(rdProc138North),
	.empty(emptyProc138North),
	.dataOut(dataInProc138North));

	//FIFO 139 TO 138 
fifo fifo_proc139_to_proc138(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc139West),
	.full(fullProc139West),
	.dataIn(dataOutProc139West),
	.rd(rdProc138East),
	.empty(emptyProc138East),
	.dataOut(dataInProc138East));
	
	//FIFO 138 TO 139
fifo fifo_proc138_to_proc139(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc138East),
	.full(fullProc138East),
	.dataIn(dataOutProc138East),
	.rd(rdProc139West),
	.empty(emptyProc139West),
	.dataOut(dataInProc139West));
	
	//FIFO 139 TO 126 
fifo fifo_proc139_to_proc126(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc139North),
	.full(fullProc139North),
	.dataIn(dataOutProc139North),
	.rd(rdProc126South),
	.empty(emptyProc126South),
	.dataOut(dataInProc126South));
	
	//FIFO 126 TO 139
fifo fifo_proc126_to_proc139(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc126South),
	.full(fullProc126South),
	.dataIn(dataOutProc126South),
	.rd(rdProc139North),
	.empty(emptyProc139North),
	.dataOut(dataInProc139North));

	//FIFO 140 TO 139 
fifo fifo_proc140_to_proc139(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc140West),
	.full(fullProc140West),
	.dataIn(dataOutProc140West),
	.rd(rdProc139East),
	.empty(emptyProc139East),
	.dataOut(dataInProc139East));
	
	//FIFO 139 TO 140
fifo fifo_proc139_to_proc140(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc139East),
	.full(fullProc139East),
	.dataIn(dataOutProc139East),
	.rd(rdProc140West),
	.empty(emptyProc140West),
	.dataOut(dataInProc140West));
	
	//FIFO 140 TO 127 
fifo fifo_proc140_to_proc127(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc140North),
	.full(fullProc140North),
	.dataIn(dataOutProc140North),
	.rd(rdProc127South),
	.empty(emptyProc127South),
	.dataOut(dataInProc127South));
	
	//FIFO 127 TO 140
fifo fifo_proc127_to_proc140(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc127South),
	.full(fullProc127South),
	.dataIn(dataOutProc127South),
	.rd(rdProc140North),
	.empty(emptyProc140North),
	.dataOut(dataInProc140North));

	//FIFO 141 TO 140 
fifo fifo_proc141_to_proc140(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc141West),
	.full(fullProc141West),
	.dataIn(dataOutProc141West),
	.rd(rdProc140East),
	.empty(emptyProc140East),
	.dataOut(dataInProc140East));
	
	//FIFO 140 TO 141
fifo fifo_proc140_to_proc141(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc140East),
	.full(fullProc140East),
	.dataIn(dataOutProc140East),
	.rd(rdProc141West),
	.empty(emptyProc141West),
	.dataOut(dataInProc141West));
	
	//FIFO 141 TO 128 
fifo fifo_proc141_to_proc128(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc141North),
	.full(fullProc141North),
	.dataIn(dataOutProc141North),
	.rd(rdProc128South),
	.empty(emptyProc128South),
	.dataOut(dataInProc128South));
	
	//FIFO 128 TO 141
fifo fifo_proc128_to_proc141(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc128South),
	.full(fullProc128South),
	.dataIn(dataOutProc128South),
	.rd(rdProc141North),
	.empty(emptyProc141North),
	.dataOut(dataInProc141North));

	//FIFO 142 TO 141 
fifo fifo_proc142_to_proc141(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc142West),
	.full(fullProc142West),
	.dataIn(dataOutProc142West),
	.rd(rdProc141East),
	.empty(emptyProc141East),
	.dataOut(dataInProc141East));
	
	//FIFO 141 TO 142
fifo fifo_proc141_to_proc142(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc141East),
	.full(fullProc141East),
	.dataIn(dataOutProc141East),
	.rd(rdProc142West),
	.empty(emptyProc142West),
	.dataOut(dataInProc142West));
	
	//FIFO 142 TO 129 
fifo fifo_proc142_to_proc129(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc142North),
	.full(fullProc142North),
	.dataIn(dataOutProc142North),
	.rd(rdProc129South),
	.empty(emptyProc129South),
	.dataOut(dataInProc129South));
	
	//FIFO 129 TO 142
fifo fifo_proc129_to_proc142(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc129South),
	.full(fullProc129South),
	.dataIn(dataOutProc129South),
	.rd(rdProc142North),
	.empty(emptyProc142North),
	.dataOut(dataInProc142North));

	//FIFO 143 TO 130 
fifo fifo_proc143_to_proc130(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc143North),
	.full(fullProc143North),
	.dataIn(dataOutProc143North),
	.rd(rdProc130South),
	.empty(emptyProc130South),
	.dataOut(dataInProc130South));
	
	//FIFO 130 TO 143
fifo fifo_proc130_to_proc143(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc130South),
	.full(fullProc130South),
	.dataIn(dataOutProc130South),
	.rd(rdProc143North),
	.empty(emptyProc143North),
	.dataOut(dataInProc143North));

	//FIFO 144 TO 143 
fifo fifo_proc144_to_proc143(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc144West),
	.full(fullProc144West),
	.dataIn(dataOutProc144West),
	.rd(rdProc143East),
	.empty(emptyProc143East),
	.dataOut(dataInProc143East));
	
	//FIFO 143 TO 144
fifo fifo_proc143_to_proc144(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc143East),
	.full(fullProc143East),
	.dataIn(dataOutProc143East),
	.rd(rdProc144West),
	.empty(emptyProc144West),
	.dataOut(dataInProc144West));
	
	//FIFO 144 TO 131 
fifo fifo_proc144_to_proc131(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc144North),
	.full(fullProc144North),
	.dataIn(dataOutProc144North),
	.rd(rdProc131South),
	.empty(emptyProc131South),
	.dataOut(dataInProc131South));
	
	//FIFO 131 TO 144
fifo fifo_proc131_to_proc144(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc131South),
	.full(fullProc131South),
	.dataIn(dataOutProc131South),
	.rd(rdProc144North),
	.empty(emptyProc144North),
	.dataOut(dataInProc144North));

	//FIFO 145 TO 144 
fifo fifo_proc145_to_proc144(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc145West),
	.full(fullProc145West),
	.dataIn(dataOutProc145West),
	.rd(rdProc144East),
	.empty(emptyProc144East),
	.dataOut(dataInProc144East));
	
	//FIFO 144 TO 145
fifo fifo_proc144_to_proc145(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc144East),
	.full(fullProc144East),
	.dataIn(dataOutProc144East),
	.rd(rdProc145West),
	.empty(emptyProc145West),
	.dataOut(dataInProc145West));
	
	//FIFO 145 TO 132 
fifo fifo_proc145_to_proc132(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc145North),
	.full(fullProc145North),
	.dataIn(dataOutProc145North),
	.rd(rdProc132South),
	.empty(emptyProc132South),
	.dataOut(dataInProc132South));
	
	//FIFO 132 TO 145
fifo fifo_proc132_to_proc145(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc132South),
	.full(fullProc132South),
	.dataIn(dataOutProc132South),
	.rd(rdProc145North),
	.empty(emptyProc145North),
	.dataOut(dataInProc145North));

	//FIFO 146 TO 145 
fifo fifo_proc146_to_proc145(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc146West),
	.full(fullProc146West),
	.dataIn(dataOutProc146West),
	.rd(rdProc145East),
	.empty(emptyProc145East),
	.dataOut(dataInProc145East));
	
	//FIFO 145 TO 146
fifo fifo_proc145_to_proc146(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc145East),
	.full(fullProc145East),
	.dataIn(dataOutProc145East),
	.rd(rdProc146West),
	.empty(emptyProc146West),
	.dataOut(dataInProc146West));
	
	//FIFO 146 TO 133 
fifo fifo_proc146_to_proc133(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc146North),
	.full(fullProc146North),
	.dataIn(dataOutProc146North),
	.rd(rdProc133South),
	.empty(emptyProc133South),
	.dataOut(dataInProc133South));
	
	//FIFO 133 TO 146
fifo fifo_proc133_to_proc146(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc133South),
	.full(fullProc133South),
	.dataIn(dataOutProc133South),
	.rd(rdProc146North),
	.empty(emptyProc146North),
	.dataOut(dataInProc146North));

	//FIFO 147 TO 146 
fifo fifo_proc147_to_proc146(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc147West),
	.full(fullProc147West),
	.dataIn(dataOutProc147West),
	.rd(rdProc146East),
	.empty(emptyProc146East),
	.dataOut(dataInProc146East));
	
	//FIFO 146 TO 147
fifo fifo_proc146_to_proc147(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc146East),
	.full(fullProc146East),
	.dataIn(dataOutProc146East),
	.rd(rdProc147West),
	.empty(emptyProc147West),
	.dataOut(dataInProc147West));
	
	//FIFO 147 TO 134 
fifo fifo_proc147_to_proc134(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc147North),
	.full(fullProc147North),
	.dataIn(dataOutProc147North),
	.rd(rdProc134South),
	.empty(emptyProc134South),
	.dataOut(dataInProc134South));
	
	//FIFO 134 TO 147
fifo fifo_proc134_to_proc147(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc134South),
	.full(fullProc134South),
	.dataIn(dataOutProc134South),
	.rd(rdProc147North),
	.empty(emptyProc147North),
	.dataOut(dataInProc147North));

	//FIFO 148 TO 147 
fifo fifo_proc148_to_proc147(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc148West),
	.full(fullProc148West),
	.dataIn(dataOutProc148West),
	.rd(rdProc147East),
	.empty(emptyProc147East),
	.dataOut(dataInProc147East));
	
	//FIFO 147 TO 148
fifo fifo_proc147_to_proc148(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc147East),
	.full(fullProc147East),
	.dataIn(dataOutProc147East),
	.rd(rdProc148West),
	.empty(emptyProc148West),
	.dataOut(dataInProc148West));
	
	//FIFO 148 TO 135 
fifo fifo_proc148_to_proc135(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc148North),
	.full(fullProc148North),
	.dataIn(dataOutProc148North),
	.rd(rdProc135South),
	.empty(emptyProc135South),
	.dataOut(dataInProc135South));
	
	//FIFO 135 TO 148
fifo fifo_proc135_to_proc148(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc135South),
	.full(fullProc135South),
	.dataIn(dataOutProc135South),
	.rd(rdProc148North),
	.empty(emptyProc148North),
	.dataOut(dataInProc148North));

	//FIFO 149 TO 148 
fifo fifo_proc149_to_proc148(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc149West),
	.full(fullProc149West),
	.dataIn(dataOutProc149West),
	.rd(rdProc148East),
	.empty(emptyProc148East),
	.dataOut(dataInProc148East));
	
	//FIFO 148 TO 149
fifo fifo_proc148_to_proc149(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc148East),
	.full(fullProc148East),
	.dataIn(dataOutProc148East),
	.rd(rdProc149West),
	.empty(emptyProc149West),
	.dataOut(dataInProc149West));
	
	//FIFO 149 TO 136 
fifo fifo_proc149_to_proc136(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc149North),
	.full(fullProc149North),
	.dataIn(dataOutProc149North),
	.rd(rdProc136South),
	.empty(emptyProc136South),
	.dataOut(dataInProc136South));
	
	//FIFO 136 TO 149
fifo fifo_proc136_to_proc149(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc136South),
	.full(fullProc136South),
	.dataIn(dataOutProc136South),
	.rd(rdProc149North),
	.empty(emptyProc149North),
	.dataOut(dataInProc149North));

	//FIFO 150 TO 149 
fifo fifo_proc150_to_proc149(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc150West),
	.full(fullProc150West),
	.dataIn(dataOutProc150West),
	.rd(rdProc149East),
	.empty(emptyProc149East),
	.dataOut(dataInProc149East));
	
	//FIFO 149 TO 150
fifo fifo_proc149_to_proc150(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc149East),
	.full(fullProc149East),
	.dataIn(dataOutProc149East),
	.rd(rdProc150West),
	.empty(emptyProc150West),
	.dataOut(dataInProc150West));
	
	//FIFO 150 TO 137 
fifo fifo_proc150_to_proc137(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc150North),
	.full(fullProc150North),
	.dataIn(dataOutProc150North),
	.rd(rdProc137South),
	.empty(emptyProc137South),
	.dataOut(dataInProc137South));
	
	//FIFO 137 TO 150
fifo fifo_proc137_to_proc150(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc137South),
	.full(fullProc137South),
	.dataIn(dataOutProc137South),
	.rd(rdProc150North),
	.empty(emptyProc150North),
	.dataOut(dataInProc150North));

	//FIFO 151 TO 150 
fifo fifo_proc151_to_proc150(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc151West),
	.full(fullProc151West),
	.dataIn(dataOutProc151West),
	.rd(rdProc150East),
	.empty(emptyProc150East),
	.dataOut(dataInProc150East));
	
	//FIFO 150 TO 151
fifo fifo_proc150_to_proc151(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc150East),
	.full(fullProc150East),
	.dataIn(dataOutProc150East),
	.rd(rdProc151West),
	.empty(emptyProc151West),
	.dataOut(dataInProc151West));
	
	//FIFO 151 TO 138 
fifo fifo_proc151_to_proc138(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc151North),
	.full(fullProc151North),
	.dataIn(dataOutProc151North),
	.rd(rdProc138South),
	.empty(emptyProc138South),
	.dataOut(dataInProc138South));
	
	//FIFO 138 TO 151
fifo fifo_proc138_to_proc151(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc138South),
	.full(fullProc138South),
	.dataIn(dataOutProc138South),
	.rd(rdProc151North),
	.empty(emptyProc151North),
	.dataOut(dataInProc151North));

	//FIFO 152 TO 151 
fifo fifo_proc152_to_proc151(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc152West),
	.full(fullProc152West),
	.dataIn(dataOutProc152West),
	.rd(rdProc151East),
	.empty(emptyProc151East),
	.dataOut(dataInProc151East));
	
	//FIFO 151 TO 152
fifo fifo_proc151_to_proc152(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc151East),
	.full(fullProc151East),
	.dataIn(dataOutProc151East),
	.rd(rdProc152West),
	.empty(emptyProc152West),
	.dataOut(dataInProc152West));
	
	//FIFO 152 TO 139 
fifo fifo_proc152_to_proc139(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc152North),
	.full(fullProc152North),
	.dataIn(dataOutProc152North),
	.rd(rdProc139South),
	.empty(emptyProc139South),
	.dataOut(dataInProc139South));
	
	//FIFO 139 TO 152
fifo fifo_proc139_to_proc152(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc139South),
	.full(fullProc139South),
	.dataIn(dataOutProc139South),
	.rd(rdProc152North),
	.empty(emptyProc152North),
	.dataOut(dataInProc152North));

	//FIFO 153 TO 152 
fifo fifo_proc153_to_proc152(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc153West),
	.full(fullProc153West),
	.dataIn(dataOutProc153West),
	.rd(rdProc152East),
	.empty(emptyProc152East),
	.dataOut(dataInProc152East));
	
	//FIFO 152 TO 153
fifo fifo_proc152_to_proc153(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc152East),
	.full(fullProc152East),
	.dataIn(dataOutProc152East),
	.rd(rdProc153West),
	.empty(emptyProc153West),
	.dataOut(dataInProc153West));
	
	//FIFO 153 TO 140 
fifo fifo_proc153_to_proc140(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc153North),
	.full(fullProc153North),
	.dataIn(dataOutProc153North),
	.rd(rdProc140South),
	.empty(emptyProc140South),
	.dataOut(dataInProc140South));
	
	//FIFO 140 TO 153
fifo fifo_proc140_to_proc153(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc140South),
	.full(fullProc140South),
	.dataIn(dataOutProc140South),
	.rd(rdProc153North),
	.empty(emptyProc153North),
	.dataOut(dataInProc153North));

	//FIFO 154 TO 153 
fifo fifo_proc154_to_proc153(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc154West),
	.full(fullProc154West),
	.dataIn(dataOutProc154West),
	.rd(rdProc153East),
	.empty(emptyProc153East),
	.dataOut(dataInProc153East));
	
	//FIFO 153 TO 154
fifo fifo_proc153_to_proc154(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc153East),
	.full(fullProc153East),
	.dataIn(dataOutProc153East),
	.rd(rdProc154West),
	.empty(emptyProc154West),
	.dataOut(dataInProc154West));
	
	//FIFO 154 TO 141 
fifo fifo_proc154_to_proc141(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc154North),
	.full(fullProc154North),
	.dataIn(dataOutProc154North),
	.rd(rdProc141South),
	.empty(emptyProc141South),
	.dataOut(dataInProc141South));
	
	//FIFO 141 TO 154
fifo fifo_proc141_to_proc154(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc141South),
	.full(fullProc141South),
	.dataIn(dataOutProc141South),
	.rd(rdProc154North),
	.empty(emptyProc154North),
	.dataOut(dataInProc154North));

	//FIFO 155 TO 154 
fifo fifo_proc155_to_proc154(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc155West),
	.full(fullProc155West),
	.dataIn(dataOutProc155West),
	.rd(rdProc154East),
	.empty(emptyProc154East),
	.dataOut(dataInProc154East));
	
	//FIFO 154 TO 155
fifo fifo_proc154_to_proc155(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc154East),
	.full(fullProc154East),
	.dataIn(dataOutProc154East),
	.rd(rdProc155West),
	.empty(emptyProc155West),
	.dataOut(dataInProc155West));
	
	//FIFO 155 TO 142 
fifo fifo_proc155_to_proc142(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc155North),
	.full(fullProc155North),
	.dataIn(dataOutProc155North),
	.rd(rdProc142South),
	.empty(emptyProc142South),
	.dataOut(dataInProc142South));
	
	//FIFO 142 TO 155
fifo fifo_proc142_to_proc155(
	.clk(clk),
	.resetn(resetn),
	.wr(wrProc142South),
	.full(fullProc142South),
	.dataIn(dataOutProc142South),
	.rd(rdProc155North),
	.empty(emptyProc155North),
	.dataOut(dataInProc155North));

	/**************** Boot loader ********************/
	/*******Boot up each processor one by one*********/
	always@(posedge clk)
	begin
	case(processor_select)
		0: begin
			boot_iwe0 = ~resetn;
			boot_dwe0 = ~resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		1: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = ~resetn;
			boot_dwe1 = ~resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		2: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = ~resetn;
			boot_dwe2 = ~resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		3: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = ~resetn;
			boot_dwe3 = ~resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		4: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = ~resetn;
			boot_dwe4 = ~resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		5: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = ~resetn;
			boot_dwe5 = ~resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		6: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = ~resetn;
			boot_dwe6 = ~resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		7: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = ~resetn;
			boot_dwe7 = ~resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		8: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = ~resetn;
			boot_dwe8 = ~resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		9: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = ~resetn;
			boot_dwe9 = ~resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		10: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = ~resetn;
			boot_dwe10 = ~resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		11: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = ~resetn;
			boot_dwe11 = ~resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		12: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = ~resetn;
			boot_dwe12 = ~resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		13: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = ~resetn;
			boot_dwe13 = ~resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		14: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = ~resetn;
			boot_dwe14 = ~resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		15: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = ~resetn;
			boot_dwe15 = ~resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		16: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = ~resetn;
			boot_dwe16 = ~resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		17: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = ~resetn;
			boot_dwe17 = ~resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		18: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = ~resetn;
			boot_dwe18 = ~resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		19: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = ~resetn;
			boot_dwe19 = ~resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		20: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = ~resetn;
			boot_dwe20 = ~resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		21: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = ~resetn;
			boot_dwe21 = ~resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		22: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = ~resetn;
			boot_dwe22 = ~resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		23: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = ~resetn;
			boot_dwe23 = ~resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		24: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = ~resetn;
			boot_dwe24 = ~resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		25: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = ~resetn;
			boot_dwe25 = ~resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		26: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = ~resetn;
			boot_dwe26 = ~resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		27: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = ~resetn;
			boot_dwe27 = ~resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		28: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = ~resetn;
			boot_dwe28 = ~resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		29: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = ~resetn;
			boot_dwe29 = ~resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		30: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = ~resetn;
			boot_dwe30 = ~resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		31: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = ~resetn;
			boot_dwe31 = ~resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		32: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = ~resetn;
			boot_dwe32 = ~resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		33: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = ~resetn;
			boot_dwe33 = ~resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		34: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = ~resetn;
			boot_dwe34 = ~resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		35: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = ~resetn;
			boot_dwe35 = ~resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		36: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = ~resetn;
			boot_dwe36 = ~resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		37: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = ~resetn;
			boot_dwe37 = ~resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		38: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = ~resetn;
			boot_dwe38 = ~resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		39: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = ~resetn;
			boot_dwe39 = ~resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		40: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = ~resetn;
			boot_dwe40 = ~resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		41: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = ~resetn;
			boot_dwe41 = ~resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		42: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = ~resetn;
			boot_dwe42 = ~resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		43: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = ~resetn;
			boot_dwe43 = ~resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		44: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = ~resetn;
			boot_dwe44 = ~resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		45: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = ~resetn;
			boot_dwe45 = ~resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		46: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = ~resetn;
			boot_dwe46 = ~resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		47: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = ~resetn;
			boot_dwe47 = ~resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		48: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = ~resetn;
			boot_dwe48 = ~resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		49: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = ~resetn;
			boot_dwe49 = ~resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		50: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = ~resetn;
			boot_dwe50 = ~resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		51: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = ~resetn;
			boot_dwe51 = ~resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		52: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = ~resetn;
			boot_dwe52 = ~resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		53: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = ~resetn;
			boot_dwe53 = ~resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		54: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = ~resetn;
			boot_dwe54 = ~resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		55: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = ~resetn;
			boot_dwe55 = ~resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		56: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = ~resetn;
			boot_dwe56 = ~resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		57: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = ~resetn;
			boot_dwe57 = ~resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		58: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = ~resetn;
			boot_dwe58 = ~resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		59: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = ~resetn;
			boot_dwe59 = ~resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		60: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = ~resetn;
			boot_dwe60 = ~resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		61: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = ~resetn;
			boot_dwe61 = ~resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		62: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = ~resetn;
			boot_dwe62 = ~resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		63: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = ~resetn;
			boot_dwe63 = ~resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		64: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = ~resetn;
			boot_dwe64 = ~resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		65: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = ~resetn;
			boot_dwe65 = ~resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		66: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = ~resetn;
			boot_dwe66 = ~resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		67: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = ~resetn;
			boot_dwe67 = ~resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		68: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = ~resetn;
			boot_dwe68 = ~resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		69: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = ~resetn;
			boot_dwe69 = ~resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		70: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = ~resetn;
			boot_dwe70 = ~resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		71: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = ~resetn;
			boot_dwe71 = ~resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		72: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = ~resetn;
			boot_dwe72 = ~resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		73: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = ~resetn;
			boot_dwe73 = ~resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		74: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = ~resetn;
			boot_dwe74 = ~resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		75: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = ~resetn;
			boot_dwe75 = ~resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		76: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = ~resetn;
			boot_dwe76 = ~resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		77: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = ~resetn;
			boot_dwe77 = ~resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		78: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = ~resetn;
			boot_dwe78 = ~resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		79: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = ~resetn;
			boot_dwe79 = ~resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		80: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = ~resetn;
			boot_dwe80 = ~resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		81: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = ~resetn;
			boot_dwe81 = ~resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		82: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = ~resetn;
			boot_dwe82 = ~resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		83: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = ~resetn;
			boot_dwe83 = ~resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		84: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = ~resetn;
			boot_dwe84 = ~resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		85: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = ~resetn;
			boot_dwe85 = ~resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		86: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = ~resetn;
			boot_dwe86 = ~resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		87: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = ~resetn;
			boot_dwe87 = ~resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		88: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = ~resetn;
			boot_dwe88 = ~resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		89: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = ~resetn;
			boot_dwe89 = ~resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		90: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = ~resetn;
			boot_dwe90 = ~resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		91: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = ~resetn;
			boot_dwe91 = ~resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		92: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = ~resetn;
			boot_dwe92 = ~resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		93: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = ~resetn;
			boot_dwe93 = ~resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		94: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = ~resetn;
			boot_dwe94 = ~resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		95: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = ~resetn;
			boot_dwe95 = ~resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		96: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = ~resetn;
			boot_dwe96 = ~resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		97: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = ~resetn;
			boot_dwe97 = ~resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		98: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = ~resetn;
			boot_dwe98 = ~resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		99: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = ~resetn;
			boot_dwe99 = ~resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		100: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = ~resetn;
			boot_dwe100 = ~resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		101: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = ~resetn;
			boot_dwe101 = ~resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		102: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = ~resetn;
			boot_dwe102 = ~resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		103: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = ~resetn;
			boot_dwe103 = ~resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		104: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = ~resetn;
			boot_dwe104 = ~resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		105: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = ~resetn;
			boot_dwe105 = ~resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		106: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = ~resetn;
			boot_dwe106 = ~resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		107: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = ~resetn;
			boot_dwe107 = ~resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		108: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = ~resetn;
			boot_dwe108 = ~resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		109: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = ~resetn;
			boot_dwe109 = ~resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		110: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = ~resetn;
			boot_dwe110 = ~resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		111: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = ~resetn;
			boot_dwe111 = ~resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		112: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = ~resetn;
			boot_dwe112 = ~resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		113: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = ~resetn;
			boot_dwe113 = ~resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		114: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = ~resetn;
			boot_dwe114 = ~resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		115: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = ~resetn;
			boot_dwe115 = ~resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		116: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = ~resetn;
			boot_dwe116 = ~resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		117: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = ~resetn;
			boot_dwe117 = ~resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		118: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = ~resetn;
			boot_dwe118 = ~resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		119: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = ~resetn;
			boot_dwe119 = ~resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		120: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = ~resetn;
			boot_dwe120 = ~resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		121: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = ~resetn;
			boot_dwe121 = ~resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		122: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = ~resetn;
			boot_dwe122 = ~resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		123: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = ~resetn;
			boot_dwe123 = ~resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		124: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = ~resetn;
			boot_dwe124 = ~resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		125: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = ~resetn;
			boot_dwe125 = ~resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		126: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = ~resetn;
			boot_dwe126 = ~resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		127: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = ~resetn;
			boot_dwe127 = ~resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		128: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = ~resetn;
			boot_dwe128 = ~resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		129: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = ~resetn;
			boot_dwe129 = ~resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		130: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = ~resetn;
			boot_dwe130 = ~resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		131: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = ~resetn;
			boot_dwe131 = ~resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		132: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = ~resetn;
			boot_dwe132 = ~resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		133: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = ~resetn;
			boot_dwe133 = ~resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		134: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = ~resetn;
			boot_dwe134 = ~resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		135: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = ~resetn;
			boot_dwe135 = ~resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		136: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = ~resetn;
			boot_dwe136 = ~resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		137: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = ~resetn;
			boot_dwe137 = ~resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		138: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = ~resetn;
			boot_dwe138 = ~resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		139: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = ~resetn;
			boot_dwe139 = ~resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		140: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = ~resetn;
			boot_dwe140 = ~resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		141: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = ~resetn;
			boot_dwe141 = ~resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		142: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = ~resetn;
			boot_dwe142 = ~resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		143: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = ~resetn;
			boot_dwe143 = ~resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		144: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = ~resetn;
			boot_dwe144 = ~resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		145: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = ~resetn;
			boot_dwe145 = ~resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		146: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = ~resetn;
			boot_dwe146 = ~resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		147: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = ~resetn;
			boot_dwe147 = ~resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		148: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = ~resetn;
			boot_dwe148 = ~resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		149: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = ~resetn;
			boot_dwe149 = ~resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		150: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = ~resetn;
			boot_dwe150 = ~resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		151: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = ~resetn;
			boot_dwe151 = ~resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		152: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = ~resetn;
			boot_dwe152 = ~resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		153: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = ~resetn;
			boot_dwe153 = ~resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		154: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = ~resetn;
			boot_dwe154 = ~resetn;
			boot_iwe155 = resetn;
			boot_dwe155 = resetn;
		end
		155: begin
			boot_iwe0 = resetn;
			boot_dwe0 = resetn;
			boot_iwe1 = resetn;
			boot_dwe1 = resetn;
			boot_iwe2 = resetn;
			boot_dwe2 = resetn;
			boot_iwe3 = resetn;
			boot_dwe3 = resetn;
			boot_iwe4 = resetn;
			boot_dwe4 = resetn;
			boot_iwe5 = resetn;
			boot_dwe5 = resetn;
			boot_iwe6 = resetn;
			boot_dwe6 = resetn;
			boot_iwe7 = resetn;
			boot_dwe7 = resetn;
			boot_iwe8 = resetn;
			boot_dwe8 = resetn;
			boot_iwe9 = resetn;
			boot_dwe9 = resetn;
			boot_iwe10 = resetn;
			boot_dwe10 = resetn;
			boot_iwe11 = resetn;
			boot_dwe11 = resetn;
			boot_iwe12 = resetn;
			boot_dwe12 = resetn;
			boot_iwe13 = resetn;
			boot_dwe13 = resetn;
			boot_iwe14 = resetn;
			boot_dwe14 = resetn;
			boot_iwe15 = resetn;
			boot_dwe15 = resetn;
			boot_iwe16 = resetn;
			boot_dwe16 = resetn;
			boot_iwe17 = resetn;
			boot_dwe17 = resetn;
			boot_iwe18 = resetn;
			boot_dwe18 = resetn;
			boot_iwe19 = resetn;
			boot_dwe19 = resetn;
			boot_iwe20 = resetn;
			boot_dwe20 = resetn;
			boot_iwe21 = resetn;
			boot_dwe21 = resetn;
			boot_iwe22 = resetn;
			boot_dwe22 = resetn;
			boot_iwe23 = resetn;
			boot_dwe23 = resetn;
			boot_iwe24 = resetn;
			boot_dwe24 = resetn;
			boot_iwe25 = resetn;
			boot_dwe25 = resetn;
			boot_iwe26 = resetn;
			boot_dwe26 = resetn;
			boot_iwe27 = resetn;
			boot_dwe27 = resetn;
			boot_iwe28 = resetn;
			boot_dwe28 = resetn;
			boot_iwe29 = resetn;
			boot_dwe29 = resetn;
			boot_iwe30 = resetn;
			boot_dwe30 = resetn;
			boot_iwe31 = resetn;
			boot_dwe31 = resetn;
			boot_iwe32 = resetn;
			boot_dwe32 = resetn;
			boot_iwe33 = resetn;
			boot_dwe33 = resetn;
			boot_iwe34 = resetn;
			boot_dwe34 = resetn;
			boot_iwe35 = resetn;
			boot_dwe35 = resetn;
			boot_iwe36 = resetn;
			boot_dwe36 = resetn;
			boot_iwe37 = resetn;
			boot_dwe37 = resetn;
			boot_iwe38 = resetn;
			boot_dwe38 = resetn;
			boot_iwe39 = resetn;
			boot_dwe39 = resetn;
			boot_iwe40 = resetn;
			boot_dwe40 = resetn;
			boot_iwe41 = resetn;
			boot_dwe41 = resetn;
			boot_iwe42 = resetn;
			boot_dwe42 = resetn;
			boot_iwe43 = resetn;
			boot_dwe43 = resetn;
			boot_iwe44 = resetn;
			boot_dwe44 = resetn;
			boot_iwe45 = resetn;
			boot_dwe45 = resetn;
			boot_iwe46 = resetn;
			boot_dwe46 = resetn;
			boot_iwe47 = resetn;
			boot_dwe47 = resetn;
			boot_iwe48 = resetn;
			boot_dwe48 = resetn;
			boot_iwe49 = resetn;
			boot_dwe49 = resetn;
			boot_iwe50 = resetn;
			boot_dwe50 = resetn;
			boot_iwe51 = resetn;
			boot_dwe51 = resetn;
			boot_iwe52 = resetn;
			boot_dwe52 = resetn;
			boot_iwe53 = resetn;
			boot_dwe53 = resetn;
			boot_iwe54 = resetn;
			boot_dwe54 = resetn;
			boot_iwe55 = resetn;
			boot_dwe55 = resetn;
			boot_iwe56 = resetn;
			boot_dwe56 = resetn;
			boot_iwe57 = resetn;
			boot_dwe57 = resetn;
			boot_iwe58 = resetn;
			boot_dwe58 = resetn;
			boot_iwe59 = resetn;
			boot_dwe59 = resetn;
			boot_iwe60 = resetn;
			boot_dwe60 = resetn;
			boot_iwe61 = resetn;
			boot_dwe61 = resetn;
			boot_iwe62 = resetn;
			boot_dwe62 = resetn;
			boot_iwe63 = resetn;
			boot_dwe63 = resetn;
			boot_iwe64 = resetn;
			boot_dwe64 = resetn;
			boot_iwe65 = resetn;
			boot_dwe65 = resetn;
			boot_iwe66 = resetn;
			boot_dwe66 = resetn;
			boot_iwe67 = resetn;
			boot_dwe67 = resetn;
			boot_iwe68 = resetn;
			boot_dwe68 = resetn;
			boot_iwe69 = resetn;
			boot_dwe69 = resetn;
			boot_iwe70 = resetn;
			boot_dwe70 = resetn;
			boot_iwe71 = resetn;
			boot_dwe71 = resetn;
			boot_iwe72 = resetn;
			boot_dwe72 = resetn;
			boot_iwe73 = resetn;
			boot_dwe73 = resetn;
			boot_iwe74 = resetn;
			boot_dwe74 = resetn;
			boot_iwe75 = resetn;
			boot_dwe75 = resetn;
			boot_iwe76 = resetn;
			boot_dwe76 = resetn;
			boot_iwe77 = resetn;
			boot_dwe77 = resetn;
			boot_iwe78 = resetn;
			boot_dwe78 = resetn;
			boot_iwe79 = resetn;
			boot_dwe79 = resetn;
			boot_iwe80 = resetn;
			boot_dwe80 = resetn;
			boot_iwe81 = resetn;
			boot_dwe81 = resetn;
			boot_iwe82 = resetn;
			boot_dwe82 = resetn;
			boot_iwe83 = resetn;
			boot_dwe83 = resetn;
			boot_iwe84 = resetn;
			boot_dwe84 = resetn;
			boot_iwe85 = resetn;
			boot_dwe85 = resetn;
			boot_iwe86 = resetn;
			boot_dwe86 = resetn;
			boot_iwe87 = resetn;
			boot_dwe87 = resetn;
			boot_iwe88 = resetn;
			boot_dwe88 = resetn;
			boot_iwe89 = resetn;
			boot_dwe89 = resetn;
			boot_iwe90 = resetn;
			boot_dwe90 = resetn;
			boot_iwe91 = resetn;
			boot_dwe91 = resetn;
			boot_iwe92 = resetn;
			boot_dwe92 = resetn;
			boot_iwe93 = resetn;
			boot_dwe93 = resetn;
			boot_iwe94 = resetn;
			boot_dwe94 = resetn;
			boot_iwe95 = resetn;
			boot_dwe95 = resetn;
			boot_iwe96 = resetn;
			boot_dwe96 = resetn;
			boot_iwe97 = resetn;
			boot_dwe97 = resetn;
			boot_iwe98 = resetn;
			boot_dwe98 = resetn;
			boot_iwe99 = resetn;
			boot_dwe99 = resetn;
			boot_iwe100 = resetn;
			boot_dwe100 = resetn;
			boot_iwe101 = resetn;
			boot_dwe101 = resetn;
			boot_iwe102 = resetn;
			boot_dwe102 = resetn;
			boot_iwe103 = resetn;
			boot_dwe103 = resetn;
			boot_iwe104 = resetn;
			boot_dwe104 = resetn;
			boot_iwe105 = resetn;
			boot_dwe105 = resetn;
			boot_iwe106 = resetn;
			boot_dwe106 = resetn;
			boot_iwe107 = resetn;
			boot_dwe107 = resetn;
			boot_iwe108 = resetn;
			boot_dwe108 = resetn;
			boot_iwe109 = resetn;
			boot_dwe109 = resetn;
			boot_iwe110 = resetn;
			boot_dwe110 = resetn;
			boot_iwe111 = resetn;
			boot_dwe111 = resetn;
			boot_iwe112 = resetn;
			boot_dwe112 = resetn;
			boot_iwe113 = resetn;
			boot_dwe113 = resetn;
			boot_iwe114 = resetn;
			boot_dwe114 = resetn;
			boot_iwe115 = resetn;
			boot_dwe115 = resetn;
			boot_iwe116 = resetn;
			boot_dwe116 = resetn;
			boot_iwe117 = resetn;
			boot_dwe117 = resetn;
			boot_iwe118 = resetn;
			boot_dwe118 = resetn;
			boot_iwe119 = resetn;
			boot_dwe119 = resetn;
			boot_iwe120 = resetn;
			boot_dwe120 = resetn;
			boot_iwe121 = resetn;
			boot_dwe121 = resetn;
			boot_iwe122 = resetn;
			boot_dwe122 = resetn;
			boot_iwe123 = resetn;
			boot_dwe123 = resetn;
			boot_iwe124 = resetn;
			boot_dwe124 = resetn;
			boot_iwe125 = resetn;
			boot_dwe125 = resetn;
			boot_iwe126 = resetn;
			boot_dwe126 = resetn;
			boot_iwe127 = resetn;
			boot_dwe127 = resetn;
			boot_iwe128 = resetn;
			boot_dwe128 = resetn;
			boot_iwe129 = resetn;
			boot_dwe129 = resetn;
			boot_iwe130 = resetn;
			boot_dwe130 = resetn;
			boot_iwe131 = resetn;
			boot_dwe131 = resetn;
			boot_iwe132 = resetn;
			boot_dwe132 = resetn;
			boot_iwe133 = resetn;
			boot_dwe133 = resetn;
			boot_iwe134 = resetn;
			boot_dwe134 = resetn;
			boot_iwe135 = resetn;
			boot_dwe135 = resetn;
			boot_iwe136 = resetn;
			boot_dwe136 = resetn;
			boot_iwe137 = resetn;
			boot_dwe137 = resetn;
			boot_iwe138 = resetn;
			boot_dwe138 = resetn;
			boot_iwe139 = resetn;
			boot_dwe139 = resetn;
			boot_iwe140 = resetn;
			boot_dwe140 = resetn;
			boot_iwe141 = resetn;
			boot_dwe141 = resetn;
			boot_iwe142 = resetn;
			boot_dwe142 = resetn;
			boot_iwe143 = resetn;
			boot_dwe143 = resetn;
			boot_iwe144 = resetn;
			boot_dwe144 = resetn;
			boot_iwe145 = resetn;
			boot_dwe145 = resetn;
			boot_iwe146 = resetn;
			boot_dwe146 = resetn;
			boot_iwe147 = resetn;
			boot_dwe147 = resetn;
			boot_iwe148 = resetn;
			boot_dwe148 = resetn;
			boot_iwe149 = resetn;
			boot_dwe149 = resetn;
			boot_iwe150 = resetn;
			boot_dwe150 = resetn;
			boot_iwe151 = resetn;
			boot_dwe151 = resetn;
			boot_iwe152 = resetn;
			boot_dwe152 = resetn;
			boot_iwe153 = resetn;
			boot_dwe153 = resetn;
			boot_iwe154 = resetn;
			boot_dwe154 = resetn;
			boot_iwe155 = ~resetn;
			boot_dwe155 = ~resetn;
		end
		156: begin
			boot_iwe0 = 0;
			boot_dwe0 = 0;
			boot_iwe1 = 0;
			boot_dwe1 = 0;
			boot_iwe2 = 0;
			boot_dwe2 = 0;
			boot_iwe3 = 0;
			boot_dwe3 = 0;
			boot_iwe4 = 0;
			boot_dwe4 = 0;
			boot_iwe5 = 0;
			boot_dwe5 = 0;
			boot_iwe6 = 0;
			boot_dwe6 = 0;
			boot_iwe7 = 0;
			boot_dwe7 = 0;
			boot_iwe8 = 0;
			boot_dwe8 = 0;
			boot_iwe9 = 0;
			boot_dwe9 = 0;
			boot_iwe10 = 0;
			boot_dwe10 = 0;
			boot_iwe11 = 0;
			boot_dwe11 = 0;
			boot_iwe12 = 0;
			boot_dwe12 = 0;
			boot_iwe13 = 0;
			boot_dwe13 = 0;
			boot_iwe14 = 0;
			boot_dwe14 = 0;
			boot_iwe15 = 0;
			boot_dwe15 = 0;
			boot_iwe16 = 0;
			boot_dwe16 = 0;
			boot_iwe17 = 0;
			boot_dwe17 = 0;
			boot_iwe18 = 0;
			boot_dwe18 = 0;
			boot_iwe19 = 0;
			boot_dwe19 = 0;
			boot_iwe20 = 0;
			boot_dwe20 = 0;
			boot_iwe21 = 0;
			boot_dwe21 = 0;
			boot_iwe22 = 0;
			boot_dwe22 = 0;
			boot_iwe23 = 0;
			boot_dwe23 = 0;
			boot_iwe24 = 0;
			boot_dwe24 = 0;
			boot_iwe25 = 0;
			boot_dwe25 = 0;
			boot_iwe26 = 0;
			boot_dwe26 = 0;
			boot_iwe27 = 0;
			boot_dwe27 = 0;
			boot_iwe28 = 0;
			boot_dwe28 = 0;
			boot_iwe29 = 0;
			boot_dwe29 = 0;
			boot_iwe30 = 0;
			boot_dwe30 = 0;
			boot_iwe31 = 0;
			boot_dwe31 = 0;
			boot_iwe32 = 0;
			boot_dwe32 = 0;
			boot_iwe33 = 0;
			boot_dwe33 = 0;
			boot_iwe34 = 0;
			boot_dwe34 = 0;
			boot_iwe35 = 0;
			boot_dwe35 = 0;
			boot_iwe36 = 0;
			boot_dwe36 = 0;
			boot_iwe37 = 0;
			boot_dwe37 = 0;
			boot_iwe38 = 0;
			boot_dwe38 = 0;
			boot_iwe39 = 0;
			boot_dwe39 = 0;
			boot_iwe40 = 0;
			boot_dwe40 = 0;
			boot_iwe41 = 0;
			boot_dwe41 = 0;
			boot_iwe42 = 0;
			boot_dwe42 = 0;
			boot_iwe43 = 0;
			boot_dwe43 = 0;
			boot_iwe44 = 0;
			boot_dwe44 = 0;
			boot_iwe45 = 0;
			boot_dwe45 = 0;
			boot_iwe46 = 0;
			boot_dwe46 = 0;
			boot_iwe47 = 0;
			boot_dwe47 = 0;
			boot_iwe48 = 0;
			boot_dwe48 = 0;
			boot_iwe49 = 0;
			boot_dwe49 = 0;
			boot_iwe50 = 0;
			boot_dwe50 = 0;
			boot_iwe51 = 0;
			boot_dwe51 = 0;
			boot_iwe52 = 0;
			boot_dwe52 = 0;
			boot_iwe53 = 0;
			boot_dwe53 = 0;
			boot_iwe54 = 0;
			boot_dwe54 = 0;
			boot_iwe55 = 0;
			boot_dwe55 = 0;
			boot_iwe56 = 0;
			boot_dwe56 = 0;
			boot_iwe57 = 0;
			boot_dwe57 = 0;
			boot_iwe58 = 0;
			boot_dwe58 = 0;
			boot_iwe59 = 0;
			boot_dwe59 = 0;
			boot_iwe60 = 0;
			boot_dwe60 = 0;
			boot_iwe61 = 0;
			boot_dwe61 = 0;
			boot_iwe62 = 0;
			boot_dwe62 = 0;
			boot_iwe63 = 0;
			boot_dwe63 = 0;
			boot_iwe64 = 0;
			boot_dwe64 = 0;
			boot_iwe65 = 0;
			boot_dwe65 = 0;
			boot_iwe66 = 0;
			boot_dwe66 = 0;
			boot_iwe67 = 0;
			boot_dwe67 = 0;
			boot_iwe68 = 0;
			boot_dwe68 = 0;
			boot_iwe69 = 0;
			boot_dwe69 = 0;
			boot_iwe70 = 0;
			boot_dwe70 = 0;
			boot_iwe71 = 0;
			boot_dwe71 = 0;
			boot_iwe72 = 0;
			boot_dwe72 = 0;
			boot_iwe73 = 0;
			boot_dwe73 = 0;
			boot_iwe74 = 0;
			boot_dwe74 = 0;
			boot_iwe75 = 0;
			boot_dwe75 = 0;
			boot_iwe76 = 0;
			boot_dwe76 = 0;
			boot_iwe77 = 0;
			boot_dwe77 = 0;
			boot_iwe78 = 0;
			boot_dwe78 = 0;
			boot_iwe79 = 0;
			boot_dwe79 = 0;
			boot_iwe80 = 0;
			boot_dwe80 = 0;
			boot_iwe81 = 0;
			boot_dwe81 = 0;
			boot_iwe82 = 0;
			boot_dwe82 = 0;
			boot_iwe83 = 0;
			boot_dwe83 = 0;
			boot_iwe84 = 0;
			boot_dwe84 = 0;
			boot_iwe85 = 0;
			boot_dwe85 = 0;
			boot_iwe86 = 0;
			boot_dwe86 = 0;
			boot_iwe87 = 0;
			boot_dwe87 = 0;
			boot_iwe88 = 0;
			boot_dwe88 = 0;
			boot_iwe89 = 0;
			boot_dwe89 = 0;
			boot_iwe90 = 0;
			boot_dwe90 = 0;
			boot_iwe91 = 0;
			boot_dwe91 = 0;
			boot_iwe92 = 0;
			boot_dwe92 = 0;
			boot_iwe93 = 0;
			boot_dwe93 = 0;
			boot_iwe94 = 0;
			boot_dwe94 = 0;
			boot_iwe95 = 0;
			boot_dwe95 = 0;
			boot_iwe96 = 0;
			boot_dwe96 = 0;
			boot_iwe97 = 0;
			boot_dwe97 = 0;
			boot_iwe98 = 0;
			boot_dwe98 = 0;
			boot_iwe99 = 0;
			boot_dwe99 = 0;
			boot_iwe100 = 0;
			boot_dwe100 = 0;
			boot_iwe101 = 0;
			boot_dwe101 = 0;
			boot_iwe102 = 0;
			boot_dwe102 = 0;
			boot_iwe103 = 0;
			boot_dwe103 = 0;
			boot_iwe104 = 0;
			boot_dwe104 = 0;
			boot_iwe105 = 0;
			boot_dwe105 = 0;
			boot_iwe106 = 0;
			boot_dwe106 = 0;
			boot_iwe107 = 0;
			boot_dwe107 = 0;
			boot_iwe108 = 0;
			boot_dwe108 = 0;
			boot_iwe109 = 0;
			boot_dwe109 = 0;
			boot_iwe110 = 0;
			boot_dwe110 = 0;
			boot_iwe111 = 0;
			boot_dwe111 = 0;
			boot_iwe112 = 0;
			boot_dwe112 = 0;
			boot_iwe113 = 0;
			boot_dwe113 = 0;
			boot_iwe114 = 0;
			boot_dwe114 = 0;
			boot_iwe115 = 0;
			boot_dwe115 = 0;
			boot_iwe116 = 0;
			boot_dwe116 = 0;
			boot_iwe117 = 0;
			boot_dwe117 = 0;
			boot_iwe118 = 0;
			boot_dwe118 = 0;
			boot_iwe119 = 0;
			boot_dwe119 = 0;
			boot_iwe120 = 0;
			boot_dwe120 = 0;
			boot_iwe121 = 0;
			boot_dwe121 = 0;
			boot_iwe122 = 0;
			boot_dwe122 = 0;
			boot_iwe123 = 0;
			boot_dwe123 = 0;
			boot_iwe124 = 0;
			boot_dwe124 = 0;
			boot_iwe125 = 0;
			boot_dwe125 = 0;
			boot_iwe126 = 0;
			boot_dwe126 = 0;
			boot_iwe127 = 0;
			boot_dwe127 = 0;
			boot_iwe128 = 0;
			boot_dwe128 = 0;
			boot_iwe129 = 0;
			boot_dwe129 = 0;
			boot_iwe130 = 0;
			boot_dwe130 = 0;
			boot_iwe131 = 0;
			boot_dwe131 = 0;
			boot_iwe132 = 0;
			boot_dwe132 = 0;
			boot_iwe133 = 0;
			boot_dwe133 = 0;
			boot_iwe134 = 0;
			boot_dwe134 = 0;
			boot_iwe135 = 0;
			boot_dwe135 = 0;
			boot_iwe136 = 0;
			boot_dwe136 = 0;
			boot_iwe137 = 0;
			boot_dwe137 = 0;
			boot_iwe138 = 0;
			boot_dwe138 = 0;
			boot_iwe139 = 0;
			boot_dwe139 = 0;
			boot_iwe140 = 0;
			boot_dwe140 = 0;
			boot_iwe141 = 0;
			boot_dwe141 = 0;
			boot_iwe142 = 0;
			boot_dwe142 = 0;
			boot_iwe143 = 0;
			boot_dwe143 = 0;
			boot_iwe144 = 0;
			boot_dwe144 = 0;
			boot_iwe145 = 0;
			boot_dwe145 = 0;
			boot_iwe146 = 0;
			boot_dwe146 = 0;
			boot_iwe147 = 0;
			boot_dwe147 = 0;
			boot_iwe148 = 0;
			boot_dwe148 = 0;
			boot_iwe149 = 0;
			boot_dwe149 = 0;
			boot_iwe150 = 0;
			boot_dwe150 = 0;
			boot_iwe151 = 0;
			boot_dwe151 = 0;
			boot_iwe152 = 0;
			boot_dwe152 = 0;
			boot_iwe153 = 0;
			boot_dwe153 = 0;
			boot_iwe154 = 0;
			boot_dwe154 = 0;
			boot_iwe155 = 0;
			boot_dwe155 = 0;
		end		
	endcase
end
endmodule