`define MAX_CLIQUESIZEBITS 5
`define MAX_VERTSBITS 12
`define MAX_PROBSBITS 16
`define MAX_PROBS (1 << `MAX_PROBSBITS)

`define MEM_ADDRBITS 26
`define MEM_WIDTHBITS 7
`define MEM_WIDTH (1 << `MEM_WIDTHBITS)
`define MEM_PROBSBITS (`MEM_ADDRBITS - (2*`MAX_VERTSBITS - `MEM_WIDTHBITS))
`define MEM_PROBS (1 << `MAX_PROBSBITS)

`define STACK_WIDTHAD 12
`define STACK_WIDTH 12
`define CACHE_HIT_LATENCY 5
`define CACHE_DEPTHBITS 8
`define CACHE_DEPTH (1 << `CACHE_DEPTHBITS)
`define CACHE_BLOCKSIZEBITS 3
`define CACHE_BLOCKSIZE (1 << `CACHE_BLOCKSIZEBITS)
`define CACHE_NBLOCKSBITS (`CACHE_DEPTHBITS - `CACHE_BLOCKSIZEBITS)
`define CACHE_NBLOCKS (1 << `CACHE_NBLOCKSBITS)
`define CACHE_TAGSIZE (`MEM_ADDRBITS - `MEM_PROBSBITS - `CACHE_DEPTHBITS)
`define MSPV_LATENCY 2

`define N_UNITSBITS 4
`define N_UNITS (1 << `N_UNITSBITS)

